/home/tom/.xschem/simulations/tb_bandgap_cascurr_cell_sw.spice