module dac_digital_interface (en_o,
    clk_i,
    rst_ni,
    randomise_en_i,
    en_i,
    VPWR,
    VGND,
    input_binary_i,
    output_binary_o,
    output_thermometer_o);
 output en_o;
 input clk_i;
 input rst_ni;
 input randomise_en_i;
 input en_i;
 input VPWR;
 input VGND;
 input [9:0] input_binary_i;
 output [1:0] output_binary_o;
 output [255:0] output_thermometer_o;

 sky130_fd_sc_hd__nor2_8 _1615_ (.A(net7),
    .B(net6),
    .Y(_1181_));
 sky130_fd_sc_hd__clkbuf_4 _1616_ (.A(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__buf_4 _1617_ (.A(net8),
    .X(_1183_));
 sky130_fd_sc_hd__clkinv_4 _1618_ (.A(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__nand2_2 _1619_ (.A(_1182_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__clkbuf_4 _1620_ (.A(net7),
    .X(_1186_));
 sky130_fd_sc_hd__buf_2 _1621_ (.A(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__buf_2 _1622_ (.A(net6),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_4 _1623_ (.A(_1183_),
    .X(_1189_));
 sky130_fd_sc_hd__o21ai_4 _1624_ (.A1(_1187_),
    .A2(_1188_),
    .B1(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__o31ai_4 _1625_ (.A1(_1186_),
    .A2(net6),
    .A3(_1183_),
    .B1(net9),
    .Y(_1191_));
 sky130_fd_sc_hd__nor2_8 _1626_ (.A(net9),
    .B(net8),
    .Y(_1192_));
 sky130_fd_sc_hd__nand2_4 _1627_ (.A(_1181_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__a22oi_4 _1628_ (.A1(_1185_),
    .A2(_1190_),
    .B1(_1191_),
    .B2(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__inv_2 _1629_ (.A(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nor2_1 _1630_ (.A(net9),
    .B(net10),
    .Y(_1196_));
 sky130_fd_sc_hd__nand3_1 _1631_ (.A(_1181_),
    .B(_1196_),
    .C(_1184_),
    .Y(_1197_));
 sky130_fd_sc_hd__buf_2 _1632_ (.A(net11),
    .X(_1198_));
 sky130_fd_sc_hd__nand2_1 _1633_ (.A(_1197_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__nor2_8 _1634_ (.A(net11),
    .B(net10),
    .Y(_1200_));
 sky130_fd_sc_hd__nand3_4 _1635_ (.A(_1181_),
    .B(_1192_),
    .C(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_2 _1636_ (.A(_1199_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__clkbuf_2 _1637_ (.A(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__nand2_2 _1638_ (.A(_1193_),
    .B(net10),
    .Y(_1204_));
 sky130_fd_sc_hd__clkbuf_2 _1639_ (.A(_1197_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_2 _1640_ (.A(_1204_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__clkbuf_4 _1641_ (.A(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__nor3_4 _1642_ (.A(_1186_),
    .B(net6),
    .C(_1183_),
    .Y(_1208_));
 sky130_fd_sc_hd__buf_4 _1643_ (.A(_1196_),
    .X(_1209_));
 sky130_fd_sc_hd__nor2_4 _1644_ (.A(net11),
    .B(net12),
    .Y(_1210_));
 sky130_fd_sc_hd__nand3_1 _1645_ (.A(_1208_),
    .B(_1209_),
    .C(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__buf_2 _1646_ (.A(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__nand3_2 _1647_ (.A(_1203_),
    .B(_1207_),
    .C(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__buf_2 _1648_ (.A(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_2 _1649_ (.A(net12),
    .X(_1215_));
 sky130_fd_sc_hd__nand2_4 _1650_ (.A(_1201_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__inv_2 _1651_ (.A(net13),
    .Y(_1217_));
 sky130_fd_sc_hd__clkbuf_2 _1652_ (.A(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__nand2_4 _1653_ (.A(_1216_),
    .B(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__inv_2 _1654_ (.A(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__buf_2 _1655_ (.A(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__buf_2 _1656_ (.A(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__o21ai_1 _1657_ (.A1(_1195_),
    .A2(_1214_),
    .B1(_1222_),
    .Y(_0514_));
 sky130_fd_sc_hd__clkinv_4 _1658_ (.A(net10),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_4 _1659_ (.A(_1210_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__clkbuf_4 _1660_ (.A(_1193_),
    .X(_1225_));
 sky130_fd_sc_hd__nor2_8 _1661_ (.A(_1224_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__buf_4 _1662_ (.A(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__nand2_2 _1663_ (.A(_1182_),
    .B(_1189_),
    .Y(_1228_));
 sky130_fd_sc_hd__o21ai_4 _1664_ (.A1(_1187_),
    .A2(_1188_),
    .B1(_1184_),
    .Y(_1229_));
 sky130_fd_sc_hd__inv_2 _1665_ (.A(_1186_),
    .Y(_1230_));
 sky130_fd_sc_hd__buf_2 _1666_ (.A(_1188_),
    .X(_1231_));
 sky130_fd_sc_hd__nand2_2 _1667_ (.A(_1230_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand3_4 _1668_ (.A(_1228_),
    .B(_1229_),
    .C(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__clkinv_4 _1669_ (.A(net9),
    .Y(_1234_));
 sky130_fd_sc_hd__o31ai_4 _1670_ (.A1(_1186_),
    .A2(net6),
    .A3(_1183_),
    .B1(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__buf_2 _1671_ (.A(net9),
    .X(_1236_));
 sky130_fd_sc_hd__nand3_4 _1672_ (.A(_1182_),
    .B(_1236_),
    .C(_1184_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_8 _1673_ (.A(_1235_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__nor2_8 _1674_ (.A(_1233_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__clkbuf_4 _1675_ (.A(_1202_),
    .X(_1240_));
 sky130_fd_sc_hd__buf_1 _1676_ (.A(_1206_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_4 _1677_ (.A(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__nand3_2 _1678_ (.A(_1239_),
    .B(_1240_),
    .C(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__o21ai_1 _1679_ (.A1(_1227_),
    .A2(_1243_),
    .B1(_1222_),
    .Y(_0513_));
 sky130_fd_sc_hd__clkbuf_4 _1680_ (.A(_1181_),
    .X(_1244_));
 sky130_fd_sc_hd__and2_4 _1681_ (.A(_1187_),
    .B(_1188_),
    .X(_1245_));
 sky130_fd_sc_hd__buf_4 _1682_ (.A(_1208_),
    .X(_1246_));
 sky130_fd_sc_hd__o21a_2 _1683_ (.A1(_1187_),
    .A2(_1188_),
    .B1(_1189_),
    .X(_1247_));
 sky130_fd_sc_hd__o22a_4 _1684_ (.A1(_1244_),
    .A2(_1245_),
    .B1(_1246_),
    .B2(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__buf_4 _1685_ (.A(_1191_),
    .X(_1249_));
 sky130_fd_sc_hd__nand2_4 _1686_ (.A(_1249_),
    .B(_1193_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _1687_ (.A(_1248_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__o21ai_1 _1688_ (.A1(_1251_),
    .A2(_1214_),
    .B1(_1222_),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _1689_ (.A(net12),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_4 _1690_ (.A(_1217_),
    .B(_1252_),
    .Y(_0511_));
 sky130_fd_sc_hd__clkbuf_2 _1691_ (.A(_1219_),
    .X(_0510_));
 sky130_fd_sc_hd__nor2_8 _1692_ (.A(_0511_),
    .B(_1201_),
    .Y(_1253_));
 sky130_fd_sc_hd__a21oi_2 _1693_ (.A1(_1216_),
    .A2(_1212_),
    .B1(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__clkbuf_2 _1694_ (.A(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_4 _1695_ (.A(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_4 _1696_ (.A(_1192_),
    .X(_1257_));
 sky130_fd_sc_hd__and4_2 _1697_ (.A(_1257_),
    .B(_1230_),
    .C(_1223_),
    .D(_1231_),
    .X(_1258_));
 sky130_fd_sc_hd__clkinv_4 _1698_ (.A(_1198_),
    .Y(_1259_));
 sky130_fd_sc_hd__buf_4 _1699_ (.A(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_1258_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand2_1 _1701_ (.A(_1211_),
    .B(net13),
    .Y(_1262_));
 sky130_fd_sc_hd__inv_2 _1702_ (.A(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__buf_2 _1703_ (.A(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__buf_2 _1704_ (.A(_1264_),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _1705_ (.A1(_1256_),
    .A2(_1261_),
    .B1(_0446_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_4 _1706_ (.A(_1198_),
    .X(_1265_));
 sky130_fd_sc_hd__nor2_8 _1707_ (.A(_1245_),
    .B(_1229_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand2_4 _1708_ (.A(_1266_),
    .B(_1209_),
    .Y(_1267_));
 sky130_fd_sc_hd__nor2_8 _1709_ (.A(_1265_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__a21o_1 _1710_ (.A1(_1216_),
    .A2(_1212_),
    .B1(_1253_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_2 _1711_ (.A(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_4 _1712_ (.A(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__buf_1 _1713_ (.A(_1262_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_4 _1714_ (.A(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__buf_1 _1715_ (.A(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__o21ai_1 _1716_ (.A1(_1268_),
    .A2(_1271_),
    .B1(_1274_),
    .Y(_0508_));
 sky130_fd_sc_hd__clkinv_4 _1717_ (.A(_1209_),
    .Y(_1275_));
 sky130_fd_sc_hd__nor2_4 _1718_ (.A(_1229_),
    .B(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__nand2_2 _1719_ (.A(_1276_),
    .B(_1260_),
    .Y(_1277_));
 sky130_fd_sc_hd__a21o_1 _1720_ (.A1(_1256_),
    .A2(_1277_),
    .B1(_0446_),
    .X(_0507_));
 sky130_fd_sc_hd__buf_2 _1721_ (.A(_1235_),
    .X(_1278_));
 sky130_fd_sc_hd__buf_4 _1722_ (.A(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__nor2_8 _1723_ (.A(_1247_),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__nand2_4 _1724_ (.A(_1280_),
    .B(_1200_),
    .Y(_1281_));
 sky130_fd_sc_hd__a21o_1 _1725_ (.A1(_1256_),
    .A2(_1281_),
    .B1(_0446_),
    .X(_0506_));
 sky130_fd_sc_hd__buf_1 _1726_ (.A(_1269_),
    .X(_1282_));
 sky130_fd_sc_hd__buf_4 _1727_ (.A(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_4 _1728_ (.A(net10),
    .X(_1284_));
 sky130_fd_sc_hd__a21oi_4 _1729_ (.A1(_1244_),
    .A2(_1257_),
    .B1(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__nand3_4 _1730_ (.A(_1233_),
    .B(_1249_),
    .C(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__buf_1 _1731_ (.A(_1202_),
    .X(_1287_));
 sky130_fd_sc_hd__buf_2 _1732_ (.A(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__nor2_4 _1733_ (.A(_1286_),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__o21ai_1 _1734_ (.A1(_1283_),
    .A2(_1289_),
    .B1(_1274_),
    .Y(_0505_));
 sky130_fd_sc_hd__buf_4 _1735_ (.A(_1203_),
    .X(_1290_));
 sky130_fd_sc_hd__o22ai_4 _1736_ (.A1(_1244_),
    .A2(_1245_),
    .B1(_1246_),
    .B2(_1247_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_2 _1737_ (.A(_1291_),
    .B(_1209_),
    .Y(_1292_));
 sky130_fd_sc_hd__nor2_4 _1738_ (.A(_1290_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__o21ai_1 _1739_ (.A1(_1283_),
    .A2(_1293_),
    .B1(_1274_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_4 _1740_ (.A(_1259_),
    .B(_1223_),
    .Y(_1294_));
 sky130_fd_sc_hd__nor2_4 _1741_ (.A(_1294_),
    .B(_1279_),
    .Y(_1295_));
 sky130_fd_sc_hd__o21ai_1 _1742_ (.A1(_1295_),
    .A2(_1271_),
    .B1(_1274_),
    .Y(_0503_));
 sky130_fd_sc_hd__buf_2 _1743_ (.A(_1249_),
    .X(_1296_));
 sky130_fd_sc_hd__and3_2 _1744_ (.A(_1296_),
    .B(_1225_),
    .C(_1200_),
    .X(_1297_));
 sky130_fd_sc_hd__o21ai_1 _1745_ (.A1(_1297_),
    .A2(_1271_),
    .B1(_1274_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand2_2 _1746_ (.A(_1193_),
    .B(_1223_),
    .Y(_1298_));
 sky130_fd_sc_hd__nand3_4 _1747_ (.A(_1182_),
    .B(_1192_),
    .C(_1284_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _1748_ (.A(_1298_),
    .B(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__clkbuf_4 _1749_ (.A(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__nand3_4 _1750_ (.A(_1230_),
    .B(_1184_),
    .C(_1231_),
    .Y(_1302_));
 sky130_fd_sc_hd__nand3_4 _1751_ (.A(_1278_),
    .B(_1237_),
    .C(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand3_4 _1752_ (.A(_1301_),
    .B(_1260_),
    .C(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__a21o_1 _1753_ (.A1(_1304_),
    .A2(_1256_),
    .B1(_0446_),
    .X(_0501_));
 sky130_fd_sc_hd__a21oi_4 _1754_ (.A1(_1225_),
    .A2(_1249_),
    .B1(_1266_),
    .Y(_1305_));
 sky130_fd_sc_hd__and3_4 _1755_ (.A(_1182_),
    .B(_1192_),
    .C(_1284_),
    .X(_1306_));
 sky130_fd_sc_hd__o21ai_4 _1756_ (.A1(_1285_),
    .A2(_1306_),
    .B1(_1259_),
    .Y(_1307_));
 sky130_fd_sc_hd__nor2_8 _1757_ (.A(_1305_),
    .B(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__buf_1 _1758_ (.A(_1273_),
    .X(_1309_));
 sky130_fd_sc_hd__o21ai_1 _1759_ (.A1(_1283_),
    .A2(_1308_),
    .B1(_1309_),
    .Y(_0500_));
 sky130_fd_sc_hd__clkbuf_2 _1760_ (.A(_1229_),
    .X(_1310_));
 sky130_fd_sc_hd__nand3_4 _1761_ (.A(_1278_),
    .B(_1237_),
    .C(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__nand3_4 _1762_ (.A(_1301_),
    .B(_1260_),
    .C(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__clkbuf_4 _1763_ (.A(_1254_),
    .X(_1313_));
 sky130_fd_sc_hd__buf_2 _1764_ (.A(_1263_),
    .X(_1314_));
 sky130_fd_sc_hd__a21o_1 _1765_ (.A1(_1312_),
    .A2(_1313_),
    .B1(_1314_),
    .X(_0499_));
 sky130_fd_sc_hd__buf_4 _1766_ (.A(_1194_),
    .X(_1315_));
 sky130_fd_sc_hd__nor2_8 _1767_ (.A(_1294_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__o21ai_1 _1768_ (.A1(_1316_),
    .A2(_1271_),
    .B1(_1309_),
    .Y(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _1769_ (.A(_1282_),
    .X(_1317_));
 sky130_fd_sc_hd__nor2_8 _1770_ (.A(_1239_),
    .B(_1307_),
    .Y(_1318_));
 sky130_fd_sc_hd__o21ai_1 _1771_ (.A1(_1317_),
    .A2(_1318_),
    .B1(_1309_),
    .Y(_0497_));
 sky130_fd_sc_hd__buf_2 _1772_ (.A(_1218_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_4 _1773_ (.A(_1250_),
    .X(_1320_));
 sky130_fd_sc_hd__a21oi_4 _1774_ (.A1(_1320_),
    .A2(_1248_),
    .B1(_1307_),
    .Y(_1321_));
 sky130_fd_sc_hd__o22ai_1 _1775_ (.A1(_1319_),
    .A2(_1226_),
    .B1(_1270_),
    .B2(_1321_),
    .Y(_0496_));
 sky130_fd_sc_hd__clkbuf_2 _1776_ (.A(_1218_),
    .X(_1322_));
 sky130_fd_sc_hd__o21ai_2 _1777_ (.A1(_1252_),
    .A2(_1200_),
    .B1(_1322_),
    .Y(_0495_));
 sky130_fd_sc_hd__a21o_1 _1778_ (.A1(_1256_),
    .A2(_1307_),
    .B1(_1314_),
    .X(_0494_));
 sky130_fd_sc_hd__and3_2 _1779_ (.A(_1257_),
    .B(_1230_),
    .C(_1231_),
    .X(_1323_));
 sky130_fd_sc_hd__inv_2 _1780_ (.A(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__clkbuf_4 _1781_ (.A(_1241_),
    .X(_1325_));
 sky130_fd_sc_hd__a21oi_4 _1782_ (.A1(_1324_),
    .A2(_1325_),
    .B1(_1290_),
    .Y(_1326_));
 sky130_fd_sc_hd__o21ai_1 _1783_ (.A1(_1317_),
    .A2(_1326_),
    .B1(_1309_),
    .Y(_0493_));
 sky130_fd_sc_hd__nor2_2 _1784_ (.A(_1236_),
    .B(_1294_),
    .Y(_1327_));
 sky130_fd_sc_hd__a21oi_4 _1785_ (.A1(_1246_),
    .A2(_1209_),
    .B1(_1259_),
    .Y(_1328_));
 sky130_fd_sc_hd__a21oi_4 _1786_ (.A1(_1327_),
    .A2(_1246_),
    .B1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__nor2_4 _1787_ (.A(_1189_),
    .B(_1244_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_2 _1788_ (.A(_1187_),
    .B(_1231_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand3_4 _1789_ (.A(_1330_),
    .B(_1234_),
    .C(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__nand3_4 _1790_ (.A(_1332_),
    .B(_1298_),
    .C(_1299_),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _1791_ (.A(_1329_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__a21o_1 _1792_ (.A1(_1334_),
    .A2(_1313_),
    .B1(_1314_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_2 _1793_ (.A(_1330_),
    .B(_1234_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand3_4 _1794_ (.A(_1335_),
    .B(_1298_),
    .C(_1299_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2_1 _1795_ (.A(_1329_),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__a21o_1 _1796_ (.A1(_1337_),
    .A2(_1313_),
    .B1(_1314_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _1797_ (.A(_1241_),
    .X(_1338_));
 sky130_fd_sc_hd__a21o_2 _1798_ (.A1(_1228_),
    .A2(_1310_),
    .B1(_1236_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_4 _1799_ (.A(_1203_),
    .X(_1340_));
 sky130_fd_sc_hd__a21oi_4 _1800_ (.A1(_1338_),
    .A2(_1339_),
    .B1(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__o21ai_1 _1801_ (.A1(_1317_),
    .A2(_1341_),
    .B1(_1309_),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_8 _1802_ (.A(_1233_),
    .B(_1249_),
    .Y(_1342_));
 sky130_fd_sc_hd__a21oi_4 _1803_ (.A1(_1342_),
    .A2(_1325_),
    .B1(_1340_),
    .Y(_1343_));
 sky130_fd_sc_hd__clkbuf_2 _1804_ (.A(_1273_),
    .X(_1344_));
 sky130_fd_sc_hd__o21ai_1 _1805_ (.A1(_1317_),
    .A2(_1343_),
    .B1(_1344_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_4 _1806_ (.A(_1291_),
    .B(_1234_),
    .Y(_1345_));
 sky130_fd_sc_hd__a21oi_2 _1807_ (.A1(_1345_),
    .A2(_1325_),
    .B1(_1340_),
    .Y(_1346_));
 sky130_fd_sc_hd__o21ai_1 _1808_ (.A1(_1317_),
    .A2(_1346_),
    .B1(_1344_),
    .Y(_0488_));
 sky130_fd_sc_hd__clkbuf_2 _1809_ (.A(_1282_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_4 _1810_ (.A(_1241_),
    .X(_1348_));
 sky130_fd_sc_hd__a21oi_2 _1811_ (.A1(_1348_),
    .A2(_1279_),
    .B1(_1290_),
    .Y(_1349_));
 sky130_fd_sc_hd__o21ai_1 _1812_ (.A1(_1347_),
    .A2(_1349_),
    .B1(_1344_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21oi_2 _1813_ (.A1(_1348_),
    .A2(_1320_),
    .B1(_1265_),
    .Y(_1350_));
 sky130_fd_sc_hd__o21ai_1 _1814_ (.A1(_1347_),
    .A2(_1350_),
    .B1(_1344_),
    .Y(_0486_));
 sky130_fd_sc_hd__and3_2 _1815_ (.A(_1278_),
    .B(_1237_),
    .C(_1302_),
    .X(_1351_));
 sky130_fd_sc_hd__a21oi_2 _1816_ (.A1(_1351_),
    .A2(_1325_),
    .B1(_1340_),
    .Y(_1352_));
 sky130_fd_sc_hd__o21ai_1 _1817_ (.A1(_1347_),
    .A2(_1352_),
    .B1(_1344_),
    .Y(_0485_));
 sky130_fd_sc_hd__clkbuf_4 _1818_ (.A(_1206_),
    .X(_1353_));
 sky130_fd_sc_hd__a21oi_2 _1819_ (.A1(_1305_),
    .A2(_1353_),
    .B1(_1340_),
    .Y(_1354_));
 sky130_fd_sc_hd__clkbuf_2 _1820_ (.A(_1273_),
    .X(_1355_));
 sky130_fd_sc_hd__o21ai_1 _1821_ (.A1(_1347_),
    .A2(_1354_),
    .B1(_1355_),
    .Y(_0484_));
 sky130_fd_sc_hd__and3_1 _1822_ (.A(_1278_),
    .B(_1237_),
    .C(_1310_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_4 _1823_ (.A(_1203_),
    .X(_1357_));
 sky130_fd_sc_hd__a21oi_2 _1824_ (.A1(_1356_),
    .A2(_1353_),
    .B1(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__o21ai_1 _1825_ (.A1(_1347_),
    .A2(_1358_),
    .B1(_1355_),
    .Y(_0483_));
 sky130_fd_sc_hd__buf_2 _1826_ (.A(_1282_),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_2 _1827_ (.A1(_1338_),
    .A2(_1315_),
    .B1(_1357_),
    .Y(_0517_));
 sky130_fd_sc_hd__o21ai_1 _1828_ (.A1(_0516_),
    .A2(_0517_),
    .B1(_1355_),
    .Y(_0482_));
 sky130_fd_sc_hd__and3_1 _1829_ (.A(_1228_),
    .B(_1310_),
    .C(_1232_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_4 _1830_ (.A(_1202_),
    .X(_0519_));
 sky130_fd_sc_hd__a31oi_2 _1831_ (.A1(_1207_),
    .A2(_0518_),
    .A3(_1250_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__o22ai_1 _1832_ (.A1(_1319_),
    .A2(_1226_),
    .B1(_1270_),
    .B2(_0520_),
    .Y(_0481_));
 sky130_fd_sc_hd__a31oi_4 _1833_ (.A1(_1207_),
    .A2(_1248_),
    .A3(_1250_),
    .B1(_0519_),
    .Y(_0521_));
 sky130_fd_sc_hd__o21ai_1 _1834_ (.A1(_0516_),
    .A2(_0521_),
    .B1(_1355_),
    .Y(_0480_));
 sky130_fd_sc_hd__clkbuf_2 _1835_ (.A(_1215_),
    .X(_0522_));
 sky130_fd_sc_hd__clkbuf_2 _1836_ (.A(net13),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_2 _1837_ (.A(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__a21o_1 _1838_ (.A1(_1265_),
    .A2(_0522_),
    .B1(_0524_),
    .X(_0479_));
 sky130_fd_sc_hd__a31o_1 _1839_ (.A1(_1205_),
    .A2(_1265_),
    .A3(_0522_),
    .B1(_0524_),
    .X(_0478_));
 sky130_fd_sc_hd__inv_2 _1840_ (.A(_1258_),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_1 _1841_ (.A(_0525_),
    .B(_1288_),
    .Y(_0526_));
 sky130_fd_sc_hd__o21ai_1 _1842_ (.A1(_0516_),
    .A2(_0526_),
    .B1(_1355_),
    .Y(_0477_));
 sky130_fd_sc_hd__clkbuf_2 _1843_ (.A(_1287_),
    .X(_0527_));
 sky130_fd_sc_hd__nand2_1 _1844_ (.A(_0527_),
    .B(_1267_),
    .Y(_0528_));
 sky130_fd_sc_hd__buf_1 _1845_ (.A(_1273_),
    .X(_0529_));
 sky130_fd_sc_hd__o21ai_1 _1846_ (.A1(_0528_),
    .A2(_1271_),
    .B1(_0529_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _1847_ (.A(_1276_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1848_ (.A(_0530_),
    .B(_1288_),
    .Y(_0531_));
 sky130_fd_sc_hd__o21ai_1 _1849_ (.A1(_0516_),
    .A2(_0531_),
    .B1(_0529_),
    .Y(_0475_));
 sky130_fd_sc_hd__nor2_4 _1850_ (.A(_1246_),
    .B(_1275_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_4 _1851_ (.A(_0532_),
    .B(_1190_),
    .Y(_0533_));
 sky130_fd_sc_hd__clkbuf_4 _1852_ (.A(_1203_),
    .X(_0534_));
 sky130_fd_sc_hd__nand2_1 _1853_ (.A(_0533_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_1 _1854_ (.A1(_0516_),
    .A2(_0535_),
    .B1(_0529_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _1855_ (.A(_1288_),
    .B(_1286_),
    .Y(_0536_));
 sky130_fd_sc_hd__clkbuf_4 _1856_ (.A(_1270_),
    .X(_0537_));
 sky130_fd_sc_hd__o21ai_1 _1857_ (.A1(_0536_),
    .A2(_0537_),
    .B1(_0529_),
    .Y(_0473_));
 sky130_fd_sc_hd__clkbuf_4 _1858_ (.A(_1282_),
    .X(_0538_));
 sky130_fd_sc_hd__nand2_1 _1859_ (.A(_1292_),
    .B(_0534_),
    .Y(_0539_));
 sky130_fd_sc_hd__o21ai_1 _1860_ (.A1(_0538_),
    .A2(_0539_),
    .B1(_0529_),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _1861_ (.A(_0532_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1862_ (.A(_0540_),
    .B(_0534_),
    .Y(_0541_));
 sky130_fd_sc_hd__clkbuf_4 _1863_ (.A(_1272_),
    .X(_0542_));
 sky130_fd_sc_hd__buf_2 _1864_ (.A(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__o21ai_1 _1865_ (.A1(_0538_),
    .A2(_0541_),
    .B1(_0543_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_1 _1866_ (.A(_1285_),
    .B(_1296_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _1867_ (.A(_1288_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__o21ai_1 _1868_ (.A1(_0545_),
    .A2(_0537_),
    .B1(_0543_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_2 _1869_ (.A(_1301_),
    .B(_1303_),
    .Y(_0546_));
 sky130_fd_sc_hd__clkbuf_2 _1870_ (.A(_1287_),
    .X(_0547_));
 sky130_fd_sc_hd__buf_2 _1871_ (.A(_1263_),
    .X(_0548_));
 sky130_fd_sc_hd__a31o_1 _1872_ (.A1(_0546_),
    .A2(_1313_),
    .A3(_0547_),
    .B1(_0548_),
    .X(_0469_));
 sky130_fd_sc_hd__o21ai_2 _1873_ (.A1(_1266_),
    .A2(_1238_),
    .B1(_1301_),
    .Y(_0549_));
 sky130_fd_sc_hd__a31o_1 _1874_ (.A1(_0549_),
    .A2(_1255_),
    .A3(_0547_),
    .B1(_0548_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_2 _1875_ (.A(_1301_),
    .B(_1311_),
    .Y(_0550_));
 sky130_fd_sc_hd__a31o_1 _1876_ (.A1(_0550_),
    .A2(_1255_),
    .A3(_0547_),
    .B1(_0548_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_2 _1877_ (.A(_1284_),
    .X(_0551_));
 sky130_fd_sc_hd__o21ai_4 _1878_ (.A1(_0551_),
    .A2(_1194_),
    .B1(_1357_),
    .Y(_0552_));
 sky130_fd_sc_hd__o21ai_1 _1879_ (.A1(_0538_),
    .A2(_0552_),
    .B1(_0543_),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_2 _1880_ (.A1(_1233_),
    .A2(_1238_),
    .B1(_1300_),
    .Y(_0553_));
 sky130_fd_sc_hd__a31o_1 _1881_ (.A1(_0553_),
    .A2(_1255_),
    .A3(_0547_),
    .B1(_1264_),
    .X(_0465_));
 sky130_fd_sc_hd__o22ai_4 _1882_ (.A1(_1285_),
    .A2(_1306_),
    .B1(_1238_),
    .B2(_1291_),
    .Y(_0554_));
 sky130_fd_sc_hd__clkbuf_2 _1883_ (.A(_1287_),
    .X(_0555_));
 sky130_fd_sc_hd__a31o_1 _1884_ (.A1(_0554_),
    .A2(_1255_),
    .A3(_0555_),
    .B1(_1264_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_2 _1885_ (.A(net13),
    .X(_0556_));
 sky130_fd_sc_hd__a31o_1 _1886_ (.A1(_1265_),
    .A2(_0551_),
    .A3(_0522_),
    .B1(_0556_),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_2 _1887_ (.A(_1259_),
    .B(_1223_),
    .Y(_0557_));
 sky130_fd_sc_hd__buf_1 _1888_ (.A(_1215_),
    .X(_0558_));
 sky130_fd_sc_hd__a31o_1 _1889_ (.A1(_0557_),
    .A2(_1225_),
    .A3(_0558_),
    .B1(_0556_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_4 _1890_ (.A(_1206_),
    .X(_0559_));
 sky130_fd_sc_hd__nand3_4 _1891_ (.A(_0534_),
    .B(_1324_),
    .C(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__o21ai_1 _1892_ (.A1(_0538_),
    .A2(_0560_),
    .B1(_0543_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand3_4 _1893_ (.A(_0534_),
    .B(_1348_),
    .C(_1332_),
    .Y(_0561_));
 sky130_fd_sc_hd__o21ai_1 _1894_ (.A1(_0561_),
    .A2(_0537_),
    .B1(_0543_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand3_4 _1895_ (.A(_0519_),
    .B(_1353_),
    .C(_1335_),
    .Y(_0562_));
 sky130_fd_sc_hd__clkbuf_2 _1896_ (.A(_0542_),
    .X(_0563_));
 sky130_fd_sc_hd__o21ai_1 _1897_ (.A1(_0562_),
    .A2(_0537_),
    .B1(_0563_),
    .Y(_0459_));
 sky130_fd_sc_hd__nand3_4 _1898_ (.A(_1290_),
    .B(_1348_),
    .C(_1339_),
    .Y(_0564_));
 sky130_fd_sc_hd__o21ai_1 _1899_ (.A1(_0564_),
    .A2(_0537_),
    .B1(_0563_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand3_4 _1900_ (.A(_0519_),
    .B(_1342_),
    .C(_1242_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21ai_1 _1901_ (.A1(_0538_),
    .A2(_0565_),
    .B1(_0563_),
    .Y(_0457_));
 sky130_fd_sc_hd__clkbuf_2 _1902_ (.A(_1269_),
    .X(_0566_));
 sky130_fd_sc_hd__nand3_4 _1903_ (.A(_1345_),
    .B(_1240_),
    .C(_1242_),
    .Y(_0567_));
 sky130_fd_sc_hd__o21ai_1 _1904_ (.A1(_0566_),
    .A2(_0567_),
    .B1(_0563_),
    .Y(_0456_));
 sky130_fd_sc_hd__clkbuf_2 _1905_ (.A(_1287_),
    .X(_0568_));
 sky130_fd_sc_hd__a41o_1 _1906_ (.A1(_1313_),
    .A2(_1279_),
    .A3(_0568_),
    .A4(_0559_),
    .B1(_1264_),
    .X(_0455_));
 sky130_fd_sc_hd__nand3_4 _1907_ (.A(_0519_),
    .B(_1353_),
    .C(_1320_),
    .Y(_0569_));
 sky130_fd_sc_hd__o21ai_1 _1908_ (.A1(_0569_),
    .A2(_1283_),
    .B1(_0563_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand3_4 _1909_ (.A(_1351_),
    .B(_1357_),
    .C(_0559_),
    .Y(_0570_));
 sky130_fd_sc_hd__clkbuf_2 _1910_ (.A(_0542_),
    .X(_0571_));
 sky130_fd_sc_hd__o21ai_1 _1911_ (.A1(_0566_),
    .A2(_0570_),
    .B1(_0571_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand3_4 _1912_ (.A(_1305_),
    .B(_1240_),
    .C(_1242_),
    .Y(_0572_));
 sky130_fd_sc_hd__o21ai_1 _1913_ (.A1(_0566_),
    .A2(_0572_),
    .B1(_0571_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand3_2 _1914_ (.A(_1356_),
    .B(_1240_),
    .C(_1242_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21ai_1 _1915_ (.A1(_0566_),
    .A2(_0573_),
    .B1(_0571_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand3_1 _1916_ (.A(_1290_),
    .B(_1348_),
    .C(_1315_),
    .Y(_0574_));
 sky130_fd_sc_hd__o21ai_1 _1917_ (.A1(_0574_),
    .A2(_1283_),
    .B1(_0571_),
    .Y(_0450_));
 sky130_fd_sc_hd__o21ai_1 _1918_ (.A1(_0566_),
    .A2(_1243_),
    .B1(_0571_),
    .Y(_0449_));
 sky130_fd_sc_hd__nor2_1 _1919_ (.A(_1238_),
    .B(_1291_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand3_2 _1920_ (.A(_0575_),
    .B(_1357_),
    .C(_0559_),
    .Y(_0576_));
 sky130_fd_sc_hd__clkbuf_2 _1921_ (.A(_0542_),
    .X(_0577_));
 sky130_fd_sc_hd__o21ai_1 _1922_ (.A1(_1270_),
    .A2(_0576_),
    .B1(_0577_),
    .Y(_0448_));
 sky130_fd_sc_hd__buf_1 _1923_ (.A(_0524_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_4 _1924_ (.A(_1216_),
    .X(_0578_));
 sky130_fd_sc_hd__inv_2 _1925_ (.A(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nor2_1 _1926_ (.A(_1261_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _1927_ (.A(_0577_),
    .B(_0580_),
    .Y(_0445_));
 sky130_fd_sc_hd__clkbuf_2 _1928_ (.A(_0578_),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_4 _1929_ (.A(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__a21oi_1 _1930_ (.A1(_1268_),
    .A2(_0582_),
    .B1(_0577_),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_2 _1931_ (.A(_1224_),
    .Y(_0583_));
 sky130_fd_sc_hd__clkbuf_2 _1932_ (.A(_1218_),
    .X(_0584_));
 sky130_fd_sc_hd__a21oi_2 _1933_ (.A1(_0583_),
    .A2(_1257_),
    .B1(_0584_),
    .Y(_0443_));
 sky130_fd_sc_hd__buf_2 _1934_ (.A(_1210_),
    .X(_0585_));
 sky130_fd_sc_hd__inv_2 _1935_ (.A(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__o21a_1 _1936_ (.A1(_0586_),
    .A2(_0533_),
    .B1(_1314_),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_1 _1937_ (.A(_1215_),
    .B(_1202_),
    .Y(_0587_));
 sky130_fd_sc_hd__clkbuf_2 _1938_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_2 _1939_ (.A(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__inv_2 _1940_ (.A(_1286_),
    .Y(_0590_));
 sky130_fd_sc_hd__a21oi_1 _1941_ (.A1(_0589_),
    .A2(_0590_),
    .B1(_0577_),
    .Y(_0441_));
 sky130_fd_sc_hd__nor2_4 _1942_ (.A(_1275_),
    .B(_1248_),
    .Y(_0591_));
 sky130_fd_sc_hd__a21oi_1 _1943_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0577_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _1944_ (.A(_1275_),
    .B(_0586_),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2_1 _1945_ (.A(_1322_),
    .B(_0592_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1946_ (.A1(_0583_),
    .A2(_1296_),
    .B1(_0584_),
    .Y(_0438_));
 sky130_fd_sc_hd__o21a_1 _1947_ (.A1(_0579_),
    .A2(_1304_),
    .B1(_0548_),
    .X(_0437_));
 sky130_fd_sc_hd__buf_2 _1948_ (.A(_0542_),
    .X(_0593_));
 sky130_fd_sc_hd__a21oi_1 _1949_ (.A1(_1308_),
    .A2(_0582_),
    .B1(_0593_),
    .Y(_0436_));
 sky130_fd_sc_hd__o21a_1 _1950_ (.A1(_0579_),
    .A2(_1312_),
    .B1(_0548_),
    .X(_0435_));
 sky130_fd_sc_hd__a21oi_1 _1951_ (.A1(_1316_),
    .A2(_0582_),
    .B1(_0593_),
    .Y(_0434_));
 sky130_fd_sc_hd__a21oi_1 _1952_ (.A1(_1318_),
    .A2(_0582_),
    .B1(_0593_),
    .Y(_0433_));
 sky130_fd_sc_hd__nor2_4 _1953_ (.A(_1198_),
    .B(_1207_),
    .Y(_0594_));
 sky130_fd_sc_hd__buf_2 _1954_ (.A(_1272_),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_2 _1955_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__a31oi_1 _1956_ (.A1(_0594_),
    .A2(_0581_),
    .A3(_1251_),
    .B1(_0596_),
    .Y(_0432_));
 sky130_fd_sc_hd__nor2_1 _1957_ (.A(_0584_),
    .B(_0583_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21oi_2 _1958_ (.A1(_1204_),
    .A2(_0585_),
    .B1(_1319_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_2 _1959_ (.A(_1324_),
    .B(_1353_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21oi_1 _1960_ (.A1(_0589_),
    .A2(_0597_),
    .B1(_0593_),
    .Y(_0429_));
 sky130_fd_sc_hd__a21oi_1 _1961_ (.A1(_0589_),
    .A2(_1333_),
    .B1(_0593_),
    .Y(_0428_));
 sky130_fd_sc_hd__buf_2 _1962_ (.A(_1272_),
    .X(_0598_));
 sky130_fd_sc_hd__buf_2 _1963_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__a21oi_1 _1964_ (.A1(_0589_),
    .A2(_1336_),
    .B1(_0599_),
    .Y(_0427_));
 sky130_fd_sc_hd__buf_2 _1965_ (.A(_0588_),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_2 _1966_ (.A(_1338_),
    .B(_1339_),
    .Y(_0601_));
 sky130_fd_sc_hd__a21oi_2 _1967_ (.A1(_0600_),
    .A2(_0601_),
    .B1(_0599_),
    .Y(_0426_));
 sky130_fd_sc_hd__clkbuf_2 _1968_ (.A(_1241_),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_2 _1969_ (.A(_1342_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__a21oi_1 _1970_ (.A1(_0600_),
    .A2(_0603_),
    .B1(_0599_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_1 _1971_ (.A(_1345_),
    .B(_0602_),
    .Y(_0604_));
 sky130_fd_sc_hd__a21oi_1 _1972_ (.A1(_0600_),
    .A2(_0604_),
    .B1(_0599_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _1973_ (.A(_1338_),
    .B(_1279_),
    .Y(_0605_));
 sky130_fd_sc_hd__a21oi_1 _1974_ (.A1(_0600_),
    .A2(_0605_),
    .B1(_0599_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _1975_ (.A(_0559_),
    .B(_1320_),
    .Y(_0606_));
 sky130_fd_sc_hd__clkbuf_2 _1976_ (.A(_0598_),
    .X(_0607_));
 sky130_fd_sc_hd__a21oi_1 _1977_ (.A1(_0606_),
    .A2(_0585_),
    .B1(_0607_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _1978_ (.A(_1351_),
    .B(_0602_),
    .Y(_0608_));
 sky130_fd_sc_hd__a21oi_1 _1979_ (.A1(_0600_),
    .A2(_0608_),
    .B1(_0607_),
    .Y(_0421_));
 sky130_fd_sc_hd__clkbuf_2 _1980_ (.A(_0588_),
    .X(_0609_));
 sky130_fd_sc_hd__nand2_1 _1981_ (.A(_1305_),
    .B(_0602_),
    .Y(_0610_));
 sky130_fd_sc_hd__a21oi_1 _1982_ (.A1(_0609_),
    .A2(_0610_),
    .B1(_0607_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _1983_ (.A(_1356_),
    .B(_0602_),
    .Y(_0611_));
 sky130_fd_sc_hd__a21oi_1 _1984_ (.A1(_0609_),
    .A2(_0611_),
    .B1(_0607_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _1985_ (.A(_1338_),
    .B(_1315_),
    .Y(_0612_));
 sky130_fd_sc_hd__a21oi_1 _1986_ (.A1(_0609_),
    .A2(_0612_),
    .B1(_0607_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _1987_ (.A(_1239_),
    .B(_1325_),
    .Y(_0613_));
 sky130_fd_sc_hd__buf_2 _1988_ (.A(_0598_),
    .X(_0614_));
 sky130_fd_sc_hd__a21oi_1 _1989_ (.A1(_0613_),
    .A2(_0609_),
    .B1(_0614_),
    .Y(_0417_));
 sky130_fd_sc_hd__nand3_2 _1990_ (.A(_1207_),
    .B(_1248_),
    .C(_1320_),
    .Y(_0615_));
 sky130_fd_sc_hd__a21oi_1 _1991_ (.A1(_0609_),
    .A2(_0615_),
    .B1(_0614_),
    .Y(_0416_));
 sky130_fd_sc_hd__nor2_1 _1992_ (.A(_0584_),
    .B(_0585_),
    .Y(_0415_));
 sky130_fd_sc_hd__a21oi_1 _1993_ (.A1(_1199_),
    .A2(_1252_),
    .B1(_1319_),
    .Y(_0414_));
 sky130_fd_sc_hd__a21oi_1 _1994_ (.A1(_0526_),
    .A2(_0582_),
    .B1(_0614_),
    .Y(_0413_));
 sky130_fd_sc_hd__clkbuf_2 _1995_ (.A(_0581_),
    .X(_0616_));
 sky130_fd_sc_hd__a21oi_1 _1996_ (.A1(_0528_),
    .A2(_0616_),
    .B1(_0614_),
    .Y(_0412_));
 sky130_fd_sc_hd__a21oi_2 _1997_ (.A1(_0531_),
    .A2(_0616_),
    .B1(_0614_),
    .Y(_0411_));
 sky130_fd_sc_hd__clkbuf_2 _1998_ (.A(_0598_),
    .X(_0617_));
 sky130_fd_sc_hd__a21oi_2 _1999_ (.A1(_0535_),
    .A2(_0616_),
    .B1(_0617_),
    .Y(_0410_));
 sky130_fd_sc_hd__a21oi_1 _2000_ (.A1(_0536_),
    .A2(_0616_),
    .B1(_0617_),
    .Y(_0409_));
 sky130_fd_sc_hd__a21oi_1 _2001_ (.A1(_0539_),
    .A2(_0616_),
    .B1(_0617_),
    .Y(_0408_));
 sky130_fd_sc_hd__clkbuf_2 _2002_ (.A(_0581_),
    .X(_0618_));
 sky130_fd_sc_hd__a21oi_1 _2003_ (.A1(_0541_),
    .A2(_0618_),
    .B1(_0617_),
    .Y(_0407_));
 sky130_fd_sc_hd__a21oi_1 _2004_ (.A1(_0545_),
    .A2(_0618_),
    .B1(_0617_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _2005_ (.A(_0546_),
    .B(_0568_),
    .Y(_0619_));
 sky130_fd_sc_hd__clkbuf_2 _2006_ (.A(_0598_),
    .X(_0620_));
 sky130_fd_sc_hd__a21oi_1 _2007_ (.A1(_0619_),
    .A2(_0618_),
    .B1(_0620_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand2_1 _2008_ (.A(_0549_),
    .B(_0527_),
    .Y(_0621_));
 sky130_fd_sc_hd__a21oi_1 _2009_ (.A1(_0621_),
    .A2(_0618_),
    .B1(_0620_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _2010_ (.A(_0550_),
    .B(_0527_),
    .Y(_0622_));
 sky130_fd_sc_hd__a21oi_1 _2011_ (.A1(_0622_),
    .A2(_0618_),
    .B1(_0620_),
    .Y(_0403_));
 sky130_fd_sc_hd__clkbuf_2 _2012_ (.A(_0578_),
    .X(_0623_));
 sky130_fd_sc_hd__a21oi_1 _2013_ (.A1(_0552_),
    .A2(_0623_),
    .B1(_0620_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _2014_ (.A(_0553_),
    .B(_0527_),
    .Y(_0624_));
 sky130_fd_sc_hd__a21oi_1 _2015_ (.A1(_0624_),
    .A2(_0623_),
    .B1(_0620_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_1 _2016_ (.A(_0554_),
    .B(_0527_),
    .Y(_0625_));
 sky130_fd_sc_hd__clkbuf_2 _2017_ (.A(_0595_),
    .X(_0626_));
 sky130_fd_sc_hd__a21oi_1 _2018_ (.A1(_0625_),
    .A2(_0623_),
    .B1(_0626_),
    .Y(_0400_));
 sky130_fd_sc_hd__o21a_1 _2019_ (.A1(_0522_),
    .A2(_0557_),
    .B1(_0524_),
    .X(_0399_));
 sky130_fd_sc_hd__nor2_1 _2020_ (.A(_1260_),
    .B(_1204_),
    .Y(_0627_));
 sky130_fd_sc_hd__o21a_1 _2021_ (.A1(_0522_),
    .A2(_0627_),
    .B1(_0524_),
    .X(_0398_));
 sky130_fd_sc_hd__a21oi_1 _2022_ (.A1(_0560_),
    .A2(_0623_),
    .B1(_0626_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_1 _2023_ (.A1(_0561_),
    .A2(_0623_),
    .B1(_0626_),
    .Y(_0396_));
 sky130_fd_sc_hd__clkbuf_2 _2024_ (.A(_0578_),
    .X(_0628_));
 sky130_fd_sc_hd__a21oi_1 _2025_ (.A1(_0562_),
    .A2(_0628_),
    .B1(_0626_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_1 _2026_ (.A1(_0564_),
    .A2(_0628_),
    .B1(_0626_),
    .Y(_0394_));
 sky130_fd_sc_hd__clkbuf_2 _2027_ (.A(_0595_),
    .X(_0629_));
 sky130_fd_sc_hd__a21oi_1 _2028_ (.A1(_0565_),
    .A2(_0628_),
    .B1(_0629_),
    .Y(_0393_));
 sky130_fd_sc_hd__a21oi_1 _2029_ (.A1(_0567_),
    .A2(_0628_),
    .B1(_0629_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _2030_ (.A(_0557_),
    .B(_1236_),
    .Y(_0630_));
 sky130_fd_sc_hd__a21oi_2 _2031_ (.A1(_0630_),
    .A2(_1252_),
    .B1(_1319_),
    .Y(_0391_));
 sky130_fd_sc_hd__a21oi_1 _2032_ (.A1(_0569_),
    .A2(_0628_),
    .B1(_0629_),
    .Y(_0390_));
 sky130_fd_sc_hd__buf_2 _2033_ (.A(_0578_),
    .X(_0631_));
 sky130_fd_sc_hd__a21oi_1 _2034_ (.A1(_0570_),
    .A2(_0631_),
    .B1(_0629_),
    .Y(_0389_));
 sky130_fd_sc_hd__a21oi_1 _2035_ (.A1(_0572_),
    .A2(_0631_),
    .B1(_0629_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_1 _2036_ (.A1(_0573_),
    .A2(_0631_),
    .B1(_0596_),
    .Y(_0387_));
 sky130_fd_sc_hd__a21oi_1 _2037_ (.A1(_0574_),
    .A2(_0631_),
    .B1(_0596_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _2038_ (.A1(_1243_),
    .A2(_0631_),
    .B1(_0596_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21oi_1 _2039_ (.A1(_0576_),
    .A2(_0581_),
    .B1(_0596_),
    .Y(_0384_));
 sky130_fd_sc_hd__nor2_1 _2040_ (.A(_0584_),
    .B(_1252_),
    .Y(_0383_));
 sky130_fd_sc_hd__nor2_8 _2041_ (.A(_1217_),
    .B(_1216_),
    .Y(_0632_));
 sky130_fd_sc_hd__clkbuf_2 _2042_ (.A(_0632_),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _2043_ (.A(_0382_),
    .B(_1261_),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _2044_ (.A(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__buf_2 _2045_ (.A(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_2 _2046_ (.A(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__nor2_1 _2047_ (.A(_1268_),
    .B(_0635_),
    .Y(_0380_));
 sky130_fd_sc_hd__and2_1 _2048_ (.A(_0382_),
    .B(_1277_),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _2049_ (.A(_1281_),
    .B(_0382_),
    .X(_0378_));
 sky130_fd_sc_hd__nor2_1 _2050_ (.A(_1289_),
    .B(_0635_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _2051_ (.A(_1293_),
    .B(_0635_),
    .Y(_0376_));
 sky130_fd_sc_hd__nor2_1 _2052_ (.A(_1295_),
    .B(_0635_),
    .Y(_0375_));
 sky130_fd_sc_hd__nor2_1 _2053_ (.A(_1297_),
    .B(_0635_),
    .Y(_0374_));
 sky130_fd_sc_hd__and2_1 _2054_ (.A(_1304_),
    .B(_0382_),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_4 _2055_ (.A(_0633_),
    .X(_0636_));
 sky130_fd_sc_hd__nor2_1 _2056_ (.A(_0636_),
    .B(_1308_),
    .Y(_0372_));
 sky130_fd_sc_hd__and2_1 _2057_ (.A(_1312_),
    .B(_0632_),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _2058_ (.A(_1316_),
    .B(_0636_),
    .Y(_0370_));
 sky130_fd_sc_hd__clkbuf_2 _2059_ (.A(_0634_),
    .X(_0637_));
 sky130_fd_sc_hd__nor2_1 _2060_ (.A(_0637_),
    .B(_1318_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _2061_ (.A(_0637_),
    .B(_1321_),
    .Y(_0368_));
 sky130_fd_sc_hd__and3_1 _2062_ (.A(_1294_),
    .B(_0556_),
    .C(_0558_),
    .X(_0367_));
 sky130_fd_sc_hd__nor2_1 _2063_ (.A(_0594_),
    .B(_0636_),
    .Y(_0366_));
 sky130_fd_sc_hd__nor2_1 _2064_ (.A(_0637_),
    .B(_1326_),
    .Y(_0365_));
 sky130_fd_sc_hd__and2_1 _2065_ (.A(_1334_),
    .B(_0632_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _2066_ (.A(_1337_),
    .B(_0632_),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_1 _2067_ (.A(_0637_),
    .B(_1341_),
    .Y(_0362_));
 sky130_fd_sc_hd__nor2_1 _2068_ (.A(_0637_),
    .B(_1343_),
    .Y(_0361_));
 sky130_fd_sc_hd__clkbuf_2 _2069_ (.A(_0634_),
    .X(_0638_));
 sky130_fd_sc_hd__nor2_1 _2070_ (.A(_0638_),
    .B(_1346_),
    .Y(_0360_));
 sky130_fd_sc_hd__nor2_1 _2071_ (.A(_1349_),
    .B(_0636_),
    .Y(_0359_));
 sky130_fd_sc_hd__nor2_1 _2072_ (.A(_1350_),
    .B(_0636_),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_0638_),
    .B(_1352_),
    .Y(_0357_));
 sky130_fd_sc_hd__nor2_1 _2074_ (.A(_0638_),
    .B(_1354_),
    .Y(_0356_));
 sky130_fd_sc_hd__nor2_1 _2075_ (.A(_0638_),
    .B(_1358_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _2076_ (.A(_0638_),
    .B(_0517_),
    .Y(_0354_));
 sky130_fd_sc_hd__nor2_1 _2077_ (.A(_0634_),
    .B(_0520_),
    .Y(_0353_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(_0634_),
    .B(_0521_),
    .Y(_0352_));
 sky130_fd_sc_hd__and3_1 _2079_ (.A(_1198_),
    .B(net13),
    .C(_1215_),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_2 _2080_ (.A(_0639_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _2081_ (.A(_1205_),
    .B(_0351_),
    .Y(_0640_));
 sky130_fd_sc_hd__inv_2 _2082_ (.A(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__clkbuf_2 _2083_ (.A(_0641_),
    .X(_0350_));
 sky130_fd_sc_hd__buf_2 _2084_ (.A(_0640_),
    .X(_0642_));
 sky130_fd_sc_hd__nor2_1 _2085_ (.A(_1258_),
    .B(_0642_),
    .Y(_0349_));
 sky130_fd_sc_hd__and3_1 _2086_ (.A(_1267_),
    .B(_1205_),
    .C(_0351_),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_1 _2087_ (.A(_0642_),
    .B(_1276_),
    .Y(_0347_));
 sky130_fd_sc_hd__and2_1 _2088_ (.A(_0350_),
    .B(_0533_),
    .X(_0346_));
 sky130_fd_sc_hd__nor2_1 _2089_ (.A(_0642_),
    .B(_0590_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _2090_ (.A(_0642_),
    .B(_0591_),
    .Y(_0344_));
 sky130_fd_sc_hd__nor2_1 _2091_ (.A(_0642_),
    .B(_0532_),
    .Y(_0343_));
 sky130_fd_sc_hd__and3_1 _2092_ (.A(_0544_),
    .B(_1205_),
    .C(_0351_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_1 _2093_ (.A(_0546_),
    .B(_0350_),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _2094_ (.A(_0549_),
    .B(_0350_),
    .X(_0340_));
 sky130_fd_sc_hd__and2_1 _2095_ (.A(_0550_),
    .B(_0641_),
    .X(_0339_));
 sky130_fd_sc_hd__o21a_1 _2096_ (.A1(_0551_),
    .A2(_1315_),
    .B1(_0350_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _2097_ (.A(_0553_),
    .B(_0641_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _2098_ (.A(_0554_),
    .B(_0641_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_4 _2099_ (.A(_0351_),
    .B(_1284_),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _2100_ (.A(_0643_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_4 _2101_ (.A(_0643_),
    .B(_1306_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _2102_ (.A(_0334_),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _2103_ (.A(_1323_),
    .B(_0644_),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _2104_ (.A(_1332_),
    .Y(_0645_));
 sky130_fd_sc_hd__nor2_1 _2105_ (.A(_0645_),
    .B(_0644_),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_1 _2106_ (.A(_1257_),
    .B(_0643_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_1 _2107_ (.A(_1280_),
    .B(_0644_),
    .Y(_0330_));
 sky130_fd_sc_hd__and2_1 _2108_ (.A(_0334_),
    .B(_1342_),
    .X(_0329_));
 sky130_fd_sc_hd__inv_2 _2109_ (.A(_1345_),
    .Y(_0646_));
 sky130_fd_sc_hd__nor2_1 _2110_ (.A(_0646_),
    .B(_0644_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _2111_ (.A(_1234_),
    .B(_0643_),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_2 _2112_ (.A(_1296_),
    .B(_0643_),
    .Y(_0326_));
 sky130_fd_sc_hd__and2_1 _2113_ (.A(_0326_),
    .B(_1302_),
    .X(_0325_));
 sky130_fd_sc_hd__o21a_1 _2114_ (.A1(_1310_),
    .A2(_1245_),
    .B1(_0326_),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_2 _2115_ (.A(_0327_),
    .B(_1189_),
    .Y(_0647_));
 sky130_fd_sc_hd__inv_2 _2116_ (.A(_0647_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor2_1 _2117_ (.A(_1244_),
    .B(_0647_),
    .Y(_0322_));
 sky130_fd_sc_hd__nor2_1 _2118_ (.A(_1230_),
    .B(_0647_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor2_1 _2119_ (.A(_1331_),
    .B(_0647_),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_1 _2120_ (.A1(_1227_),
    .A2(_0580_),
    .B1(_1322_),
    .Y(_0318_));
 sky130_fd_sc_hd__clkbuf_4 _2121_ (.A(_1253_),
    .X(_0648_));
 sky130_fd_sc_hd__a21oi_1 _2122_ (.A1(_1221_),
    .A2(_1268_),
    .B1(_0648_),
    .Y(_0317_));
 sky130_fd_sc_hd__buf_1 _2123_ (.A(_1212_),
    .X(_0649_));
 sky130_fd_sc_hd__buf_2 _2124_ (.A(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a21o_1 _2125_ (.A1(_1277_),
    .A2(_0650_),
    .B1(_0510_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_2 _2126_ (.A(_1253_),
    .X(_0651_));
 sky130_fd_sc_hd__inv_2 _2127_ (.A(_0651_),
    .Y(_0515_));
 sky130_fd_sc_hd__o31a_1 _2128_ (.A1(_0586_),
    .A2(_0533_),
    .A3(_1264_),
    .B1(_0515_),
    .X(_0315_));
 sky130_fd_sc_hd__buf_2 _2129_ (.A(_0588_),
    .X(_0652_));
 sky130_fd_sc_hd__buf_2 _2130_ (.A(_0595_),
    .X(_0653_));
 sky130_fd_sc_hd__a31oi_4 _2131_ (.A1(_0652_),
    .A2(_0590_),
    .A3(_0653_),
    .B1(_0648_),
    .Y(_0314_));
 sky130_fd_sc_hd__a31oi_1 _2132_ (.A1(_0652_),
    .A2(_0591_),
    .A3(_0653_),
    .B1(_0648_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _2133_ (.A(_0592_),
    .B(_1322_),
    .Y(_0312_));
 sky130_fd_sc_hd__or3b_2 _2134_ (.A(_0523_),
    .B(_1224_),
    .C_N(_1296_),
    .X(_0311_));
 sky130_fd_sc_hd__o31a_1 _2135_ (.A1(_0556_),
    .A2(_0579_),
    .A3(_1304_),
    .B1(_0515_),
    .X(_0310_));
 sky130_fd_sc_hd__a21oi_1 _2136_ (.A1(_1308_),
    .A2(_1221_),
    .B1(_0648_),
    .Y(_0309_));
 sky130_fd_sc_hd__o31a_1 _2137_ (.A1(_0556_),
    .A2(_0579_),
    .A3(_1312_),
    .B1(_0515_),
    .X(_0308_));
 sky130_fd_sc_hd__o21ai_1 _2138_ (.A1(_1227_),
    .A2(_1316_),
    .B1(_1222_),
    .Y(_0307_));
 sky130_fd_sc_hd__o21ai_1 _2139_ (.A1(_1227_),
    .A2(_1318_),
    .B1(_1222_),
    .Y(_0306_));
 sky130_fd_sc_hd__a31oi_1 _2140_ (.A1(_1221_),
    .A2(_0594_),
    .A3(_1251_),
    .B1(_0648_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _2141_ (.A(_0583_),
    .B(_1322_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand2_1 _2142_ (.A(_0585_),
    .B(_1218_),
    .Y(_0288_));
 sky130_fd_sc_hd__a21o_1 _2143_ (.A1(_1225_),
    .A2(_0551_),
    .B1(_0288_),
    .X(_0303_));
 sky130_fd_sc_hd__buf_1 _2144_ (.A(_0651_),
    .X(_0654_));
 sky130_fd_sc_hd__a31oi_1 _2145_ (.A1(_0652_),
    .A2(_0597_),
    .A3(_0653_),
    .B1(_0654_),
    .Y(_0302_));
 sky130_fd_sc_hd__clkbuf_2 _2146_ (.A(_1272_),
    .X(_0655_));
 sky130_fd_sc_hd__a31oi_1 _2147_ (.A1(_0652_),
    .A2(_0655_),
    .A3(_1333_),
    .B1(_0654_),
    .Y(_0301_));
 sky130_fd_sc_hd__a31oi_1 _2148_ (.A1(_0652_),
    .A2(_0655_),
    .A3(_1336_),
    .B1(_0654_),
    .Y(_0300_));
 sky130_fd_sc_hd__buf_2 _2149_ (.A(_0588_),
    .X(_0656_));
 sky130_fd_sc_hd__a31oi_1 _2150_ (.A1(_0656_),
    .A2(_0601_),
    .A3(_0653_),
    .B1(_0654_),
    .Y(_0299_));
 sky130_fd_sc_hd__a31oi_1 _2151_ (.A1(_0656_),
    .A2(_0603_),
    .A3(_0653_),
    .B1(_0654_),
    .Y(_0298_));
 sky130_fd_sc_hd__clkbuf_2 _2152_ (.A(_0595_),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_2 _2153_ (.A(_1253_),
    .X(_0658_));
 sky130_fd_sc_hd__a31oi_1 _2154_ (.A1(_0656_),
    .A2(_0604_),
    .A3(_0657_),
    .B1(_0658_),
    .Y(_0297_));
 sky130_fd_sc_hd__a31oi_1 _2155_ (.A1(_0656_),
    .A2(_0605_),
    .A3(_0657_),
    .B1(_0658_),
    .Y(_0296_));
 sky130_fd_sc_hd__a31o_1 _2156_ (.A1(_1185_),
    .A2(_1236_),
    .A3(_0551_),
    .B1(_0288_),
    .X(_0295_));
 sky130_fd_sc_hd__a31oi_1 _2157_ (.A1(_0656_),
    .A2(_0608_),
    .A3(_0657_),
    .B1(_0658_),
    .Y(_0294_));
 sky130_fd_sc_hd__clkbuf_2 _2158_ (.A(_0587_),
    .X(_0659_));
 sky130_fd_sc_hd__a31oi_1 _2159_ (.A1(_0659_),
    .A2(_0610_),
    .A3(_0657_),
    .B1(_0658_),
    .Y(_0293_));
 sky130_fd_sc_hd__a31oi_1 _2160_ (.A1(_0659_),
    .A2(_0611_),
    .A3(_0657_),
    .B1(_0658_),
    .Y(_0292_));
 sky130_fd_sc_hd__a31oi_1 _2161_ (.A1(_0659_),
    .A2(_0612_),
    .A3(_0655_),
    .B1(_0651_),
    .Y(_0291_));
 sky130_fd_sc_hd__a31oi_1 _2162_ (.A1(_0613_),
    .A2(_0659_),
    .A3(_0655_),
    .B1(_0651_),
    .Y(_0290_));
 sky130_fd_sc_hd__a31oi_1 _2163_ (.A1(_0659_),
    .A2(_0615_),
    .A3(_0655_),
    .B1(_0651_),
    .Y(_0289_));
 sky130_fd_sc_hd__or2_1 _2164_ (.A(_0511_),
    .B(_1328_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_2 _2165_ (.A(_1240_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_2 _2166_ (.A(_1212_),
    .X(_0661_));
 sky130_fd_sc_hd__a31o_1 _2167_ (.A1(_0525_),
    .A2(_0660_),
    .A3(_0661_),
    .B1(_0510_),
    .X(_0286_));
 sky130_fd_sc_hd__a31o_1 _2168_ (.A1(_0660_),
    .A2(_1267_),
    .A3(_0649_),
    .B1(_0510_),
    .X(_0285_));
 sky130_fd_sc_hd__a31o_1 _2169_ (.A1(_0530_),
    .A2(_0650_),
    .A3(_0555_),
    .B1(_0510_),
    .X(_0284_));
 sky130_fd_sc_hd__buf_1 _2170_ (.A(_1219_),
    .X(_0662_));
 sky130_fd_sc_hd__a31o_1 _2171_ (.A1(_0533_),
    .A2(_0660_),
    .A3(_0649_),
    .B1(_0662_),
    .X(_0283_));
 sky130_fd_sc_hd__a31o_1 _2172_ (.A1(_0660_),
    .A2(_1286_),
    .A3(_0649_),
    .B1(_0662_),
    .X(_0282_));
 sky130_fd_sc_hd__a31o_1 _2173_ (.A1(_1292_),
    .A2(_0547_),
    .A3(_0649_),
    .B1(_0662_),
    .X(_0281_));
 sky130_fd_sc_hd__a31o_1 _2174_ (.A1(_0540_),
    .A2(_0650_),
    .A3(_0555_),
    .B1(_0662_),
    .X(_0280_));
 sky130_fd_sc_hd__a31o_1 _2175_ (.A1(_0660_),
    .A2(_0650_),
    .A3(_0544_),
    .B1(_0662_),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_2 _2176_ (.A(_1219_),
    .X(_0663_));
 sky130_fd_sc_hd__a31o_1 _2177_ (.A1(_0546_),
    .A2(_0650_),
    .A3(_0555_),
    .B1(_0663_),
    .X(_0278_));
 sky130_fd_sc_hd__a31o_1 _2178_ (.A1(_0549_),
    .A2(_0661_),
    .A3(_0555_),
    .B1(_0663_),
    .X(_0277_));
 sky130_fd_sc_hd__a31o_1 _2179_ (.A1(_0550_),
    .A2(_0661_),
    .A3(_0568_),
    .B1(_0663_),
    .X(_0276_));
 sky130_fd_sc_hd__clkbuf_2 _2180_ (.A(_1220_),
    .X(_0664_));
 sky130_fd_sc_hd__o21ai_1 _2181_ (.A1(_1227_),
    .A2(_0552_),
    .B1(_0664_),
    .Y(_0275_));
 sky130_fd_sc_hd__a31o_1 _2182_ (.A1(_0553_),
    .A2(_0661_),
    .A3(_0568_),
    .B1(_0663_),
    .X(_0274_));
 sky130_fd_sc_hd__a31o_1 _2183_ (.A1(_0554_),
    .A2(_0661_),
    .A3(_0568_),
    .B1(_0663_),
    .X(_0273_));
 sky130_fd_sc_hd__or3_1 _2184_ (.A(_0523_),
    .B(_0558_),
    .C(_0557_),
    .X(_0272_));
 sky130_fd_sc_hd__or3_1 _2185_ (.A(_0523_),
    .B(_0558_),
    .C(_0627_),
    .X(_0271_));
 sky130_fd_sc_hd__o21ai_1 _2186_ (.A1(_1323_),
    .A2(_1214_),
    .B1(_0664_),
    .Y(_0270_));
 sky130_fd_sc_hd__o21ai_1 _2187_ (.A1(_0645_),
    .A2(_1214_),
    .B1(_0664_),
    .Y(_0269_));
 sky130_fd_sc_hd__clkbuf_2 _2188_ (.A(_1226_),
    .X(_0665_));
 sky130_fd_sc_hd__o21ai_1 _2189_ (.A1(_0665_),
    .A2(_0562_),
    .B1(_0664_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_1 _2190_ (.A1(_1280_),
    .A2(_1214_),
    .B1(_0664_),
    .Y(_0267_));
 sky130_fd_sc_hd__clkbuf_2 _2191_ (.A(_1220_),
    .X(_0666_));
 sky130_fd_sc_hd__o21ai_1 _2192_ (.A1(_0665_),
    .A2(_0565_),
    .B1(_0666_),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_1 _2193_ (.A1(_0665_),
    .A2(_0567_),
    .B1(_0666_),
    .Y(_0265_));
 sky130_fd_sc_hd__or3b_1 _2194_ (.A(_0523_),
    .B(_0558_),
    .C_N(_0630_),
    .X(_0264_));
 sky130_fd_sc_hd__o21ai_1 _2195_ (.A1(_0665_),
    .A2(_0569_),
    .B1(_0666_),
    .Y(_0263_));
 sky130_fd_sc_hd__o21ai_1 _2196_ (.A1(_1303_),
    .A2(_1213_),
    .B1(_0666_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21ai_1 _2197_ (.A1(_0665_),
    .A2(_0572_),
    .B1(_0666_),
    .Y(_0261_));
 sky130_fd_sc_hd__o21ai_1 _2198_ (.A1(_1226_),
    .A2(_0573_),
    .B1(_1221_),
    .Y(_0260_));
 sky130_fd_sc_hd__and2_1 _2199_ (.A(net2),
    .B(\lfsr_q[13] ),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(net2),
    .B(\lfsr_q[14] ),
    .X(_0002_));
 sky130_fd_sc_hd__buf_1 _2201_ (.A(\remap_control[0] ),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_4 _2202_ (.A(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__buf_2 _2203_ (.A(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_1 _2204_ (.A(\remap_control[1] ),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_4 _2205_ (.A(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__buf_2 _2206_ (.A(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_8 _2207_ (.A(_0669_),
    .B(_0672_),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _2208_ (.A(\remap_control[1] ),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_2 _2209_ (.A(_0667_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__buf_2 _2210_ (.A(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_2 _2211_ (.A(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__and2_1 _2212_ (.A(_0673_),
    .B(\remap_control[0] ),
    .X(_0677_));
 sky130_fd_sc_hd__buf_2 _2213_ (.A(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_2 _2214_ (.A(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__and3_1 _2215_ (.A(_0669_),
    .B(_0672_),
    .C(\reversed_thermometer[191] ),
    .X(_0680_));
 sky130_fd_sc_hd__a221o_1 _2216_ (.A1(\reversed_thermometer[127] ),
    .A2(_0676_),
    .B1(_0679_),
    .B2(\reversed_thermometer[63] ),
    .C1(_0680_),
    .X(_0228_));
 sky130_fd_sc_hd__and3_1 _2217_ (.A(_0669_),
    .B(_0672_),
    .C(\reversed_thermometer[190] ),
    .X(_0681_));
 sky130_fd_sc_hd__a221o_1 _2218_ (.A1(\reversed_thermometer[126] ),
    .A2(_0676_),
    .B1(_0679_),
    .B2(\reversed_thermometer[62] ),
    .C1(_0681_),
    .X(_0229_));
 sky130_fd_sc_hd__and3_1 _2219_ (.A(_0669_),
    .B(_0672_),
    .C(\reversed_thermometer[189] ),
    .X(_0682_));
 sky130_fd_sc_hd__a221o_1 _2220_ (.A1(\reversed_thermometer[125] ),
    .A2(_0676_),
    .B1(_0679_),
    .B2(\reversed_thermometer[61] ),
    .C1(_0682_),
    .X(_0230_));
 sky130_fd_sc_hd__and3_1 _2221_ (.A(_0669_),
    .B(_0672_),
    .C(\reversed_thermometer[188] ),
    .X(_0683_));
 sky130_fd_sc_hd__a221o_1 _2222_ (.A1(\reversed_thermometer[124] ),
    .A2(_0676_),
    .B1(_0679_),
    .B2(\reversed_thermometer[60] ),
    .C1(_0683_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_2 _2223_ (.A(_0668_),
    .X(_0684_));
 sky130_fd_sc_hd__buf_1 _2224_ (.A(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_2 _2225_ (.A(_0671_),
    .X(_0686_));
 sky130_fd_sc_hd__buf_1 _2226_ (.A(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__and3_1 _2227_ (.A(_0685_),
    .B(_0687_),
    .C(\reversed_thermometer[187] ),
    .X(_0688_));
 sky130_fd_sc_hd__a221o_1 _2228_ (.A1(\reversed_thermometer[123] ),
    .A2(_0676_),
    .B1(_0679_),
    .B2(\reversed_thermometer[59] ),
    .C1(_0688_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_2 _2229_ (.A(_0675_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_2 _2230_ (.A(_0678_),
    .X(_0690_));
 sky130_fd_sc_hd__and3_1 _2231_ (.A(_0685_),
    .B(_0687_),
    .C(\reversed_thermometer[186] ),
    .X(_0691_));
 sky130_fd_sc_hd__a221o_1 _2232_ (.A1(\reversed_thermometer[122] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\reversed_thermometer[58] ),
    .C1(_0691_),
    .X(_0233_));
 sky130_fd_sc_hd__and3_1 _2233_ (.A(_0685_),
    .B(_0687_),
    .C(\reversed_thermometer[185] ),
    .X(_0692_));
 sky130_fd_sc_hd__a221o_1 _2234_ (.A1(\reversed_thermometer[121] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\reversed_thermometer[57] ),
    .C1(_0692_),
    .X(_0234_));
 sky130_fd_sc_hd__and3_1 _2235_ (.A(_0685_),
    .B(_0687_),
    .C(\reversed_thermometer[184] ),
    .X(_0693_));
 sky130_fd_sc_hd__a221o_1 _2236_ (.A1(\reversed_thermometer[120] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\reversed_thermometer[56] ),
    .C1(_0693_),
    .X(_0235_));
 sky130_fd_sc_hd__and3_1 _2237_ (.A(_0685_),
    .B(_0687_),
    .C(\reversed_thermometer[183] ),
    .X(_0694_));
 sky130_fd_sc_hd__a221o_1 _2238_ (.A1(\reversed_thermometer[119] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\reversed_thermometer[55] ),
    .C1(_0694_),
    .X(_0236_));
 sky130_fd_sc_hd__buf_1 _2239_ (.A(_0684_),
    .X(_0695_));
 sky130_fd_sc_hd__buf_1 _2240_ (.A(_0686_),
    .X(_0696_));
 sky130_fd_sc_hd__and3_1 _2241_ (.A(_0695_),
    .B(_0696_),
    .C(\reversed_thermometer[182] ),
    .X(_0697_));
 sky130_fd_sc_hd__a221o_1 _2242_ (.A1(\reversed_thermometer[118] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\reversed_thermometer[54] ),
    .C1(_0697_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_2 _2243_ (.A(_0675_),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_2 _2244_ (.A(_0678_),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _2245_ (.A(_0695_),
    .B(_0696_),
    .C(\reversed_thermometer[181] ),
    .X(_0700_));
 sky130_fd_sc_hd__a221o_1 _2246_ (.A1(\reversed_thermometer[117] ),
    .A2(_0698_),
    .B1(_0699_),
    .B2(\reversed_thermometer[53] ),
    .C1(_0700_),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _2247_ (.A(_0695_),
    .B(_0696_),
    .C(\reversed_thermometer[180] ),
    .X(_0701_));
 sky130_fd_sc_hd__a221o_1 _2248_ (.A1(\reversed_thermometer[116] ),
    .A2(_0698_),
    .B1(_0699_),
    .B2(\reversed_thermometer[52] ),
    .C1(_0701_),
    .X(_0239_));
 sky130_fd_sc_hd__and3_1 _2249_ (.A(_0695_),
    .B(_0696_),
    .C(\reversed_thermometer[179] ),
    .X(_0702_));
 sky130_fd_sc_hd__a221o_1 _2250_ (.A1(\reversed_thermometer[115] ),
    .A2(_0698_),
    .B1(_0699_),
    .B2(\reversed_thermometer[51] ),
    .C1(_0702_),
    .X(_0240_));
 sky130_fd_sc_hd__and3_1 _2251_ (.A(_0695_),
    .B(_0696_),
    .C(\reversed_thermometer[178] ),
    .X(_0703_));
 sky130_fd_sc_hd__a221o_1 _2252_ (.A1(\reversed_thermometer[114] ),
    .A2(_0698_),
    .B1(_0699_),
    .B2(\reversed_thermometer[50] ),
    .C1(_0703_),
    .X(_0241_));
 sky130_fd_sc_hd__buf_1 _2253_ (.A(_0684_),
    .X(_0704_));
 sky130_fd_sc_hd__buf_1 _2254_ (.A(_0686_),
    .X(_0705_));
 sky130_fd_sc_hd__and3_1 _2255_ (.A(_0704_),
    .B(_0705_),
    .C(\reversed_thermometer[177] ),
    .X(_0706_));
 sky130_fd_sc_hd__a221o_1 _2256_ (.A1(\reversed_thermometer[113] ),
    .A2(_0698_),
    .B1(_0699_),
    .B2(\reversed_thermometer[49] ),
    .C1(_0706_),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_2 _2257_ (.A(_0675_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_2 _2258_ (.A(_0678_),
    .X(_0708_));
 sky130_fd_sc_hd__and3_1 _2259_ (.A(_0704_),
    .B(_0705_),
    .C(\reversed_thermometer[176] ),
    .X(_0709_));
 sky130_fd_sc_hd__a221o_1 _2260_ (.A1(\reversed_thermometer[112] ),
    .A2(_0707_),
    .B1(_0708_),
    .B2(\reversed_thermometer[48] ),
    .C1(_0709_),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _2261_ (.A(_0704_),
    .B(_0705_),
    .C(\reversed_thermometer[175] ),
    .X(_0710_));
 sky130_fd_sc_hd__a221o_1 _2262_ (.A1(\reversed_thermometer[111] ),
    .A2(_0707_),
    .B1(_0708_),
    .B2(\reversed_thermometer[47] ),
    .C1(_0710_),
    .X(_0244_));
 sky130_fd_sc_hd__and3_1 _2263_ (.A(_0704_),
    .B(_0705_),
    .C(\reversed_thermometer[174] ),
    .X(_0711_));
 sky130_fd_sc_hd__a221o_1 _2264_ (.A1(\reversed_thermometer[110] ),
    .A2(_0707_),
    .B1(_0708_),
    .B2(\reversed_thermometer[46] ),
    .C1(_0711_),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _2265_ (.A(_0704_),
    .B(_0705_),
    .C(\reversed_thermometer[173] ),
    .X(_0712_));
 sky130_fd_sc_hd__a221o_1 _2266_ (.A1(\reversed_thermometer[109] ),
    .A2(_0707_),
    .B1(_0708_),
    .B2(\reversed_thermometer[45] ),
    .C1(_0712_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_4 _2267_ (.A(_0668_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_1 _2268_ (.A(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_4 _2269_ (.A(_0671_),
    .X(_0715_));
 sky130_fd_sc_hd__buf_1 _2270_ (.A(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__and3_1 _2271_ (.A(_0714_),
    .B(_0716_),
    .C(\reversed_thermometer[172] ),
    .X(_0717_));
 sky130_fd_sc_hd__a221o_1 _2272_ (.A1(\reversed_thermometer[108] ),
    .A2(_0707_),
    .B1(_0708_),
    .B2(\reversed_thermometer[44] ),
    .C1(_0717_),
    .X(_0247_));
 sky130_fd_sc_hd__buf_2 _2273_ (.A(_0674_),
    .X(_0718_));
 sky130_fd_sc_hd__buf_2 _2274_ (.A(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__buf_2 _2275_ (.A(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__buf_2 _2276_ (.A(_0677_),
    .X(_0721_));
 sky130_fd_sc_hd__buf_2 _2277_ (.A(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__buf_2 _2278_ (.A(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__and3_1 _2279_ (.A(_0714_),
    .B(_0716_),
    .C(\reversed_thermometer[171] ),
    .X(_0724_));
 sky130_fd_sc_hd__a221o_1 _2280_ (.A1(\reversed_thermometer[107] ),
    .A2(_0720_),
    .B1(_0723_),
    .B2(\reversed_thermometer[43] ),
    .C1(_0724_),
    .X(_0248_));
 sky130_fd_sc_hd__and3_1 _2281_ (.A(_0714_),
    .B(_0716_),
    .C(\reversed_thermometer[170] ),
    .X(_0725_));
 sky130_fd_sc_hd__a221o_1 _2282_ (.A1(\reversed_thermometer[106] ),
    .A2(_0720_),
    .B1(_0723_),
    .B2(\reversed_thermometer[42] ),
    .C1(_0725_),
    .X(_0249_));
 sky130_fd_sc_hd__and3_1 _2283_ (.A(_0714_),
    .B(_0716_),
    .C(\reversed_thermometer[169] ),
    .X(_0726_));
 sky130_fd_sc_hd__a221o_1 _2284_ (.A1(\reversed_thermometer[105] ),
    .A2(_0720_),
    .B1(_0723_),
    .B2(\reversed_thermometer[41] ),
    .C1(_0726_),
    .X(_0250_));
 sky130_fd_sc_hd__and3_1 _2285_ (.A(_0714_),
    .B(_0716_),
    .C(\reversed_thermometer[168] ),
    .X(_0727_));
 sky130_fd_sc_hd__a221o_1 _2286_ (.A1(\reversed_thermometer[104] ),
    .A2(_0720_),
    .B1(_0723_),
    .B2(\reversed_thermometer[40] ),
    .C1(_0727_),
    .X(_0251_));
 sky130_fd_sc_hd__buf_1 _2287_ (.A(_0713_),
    .X(_0728_));
 sky130_fd_sc_hd__buf_1 _2288_ (.A(_0715_),
    .X(_0729_));
 sky130_fd_sc_hd__and3_1 _2289_ (.A(_0728_),
    .B(_0729_),
    .C(\reversed_thermometer[167] ),
    .X(_0730_));
 sky130_fd_sc_hd__a221o_1 _2290_ (.A1(\reversed_thermometer[103] ),
    .A2(_0720_),
    .B1(_0723_),
    .B2(\reversed_thermometer[39] ),
    .C1(_0730_),
    .X(_0252_));
 sky130_fd_sc_hd__buf_1 _2291_ (.A(_0719_),
    .X(_0731_));
 sky130_fd_sc_hd__buf_1 _2292_ (.A(_0722_),
    .X(_0732_));
 sky130_fd_sc_hd__and3_1 _2293_ (.A(_0728_),
    .B(_0729_),
    .C(\reversed_thermometer[166] ),
    .X(_0733_));
 sky130_fd_sc_hd__a221o_1 _2294_ (.A1(\reversed_thermometer[102] ),
    .A2(_0731_),
    .B1(_0732_),
    .B2(\reversed_thermometer[38] ),
    .C1(_0733_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _2295_ (.A(_0728_),
    .B(_0729_),
    .C(\reversed_thermometer[165] ),
    .X(_0734_));
 sky130_fd_sc_hd__a221o_1 _2296_ (.A1(\reversed_thermometer[101] ),
    .A2(_0731_),
    .B1(_0732_),
    .B2(\reversed_thermometer[37] ),
    .C1(_0734_),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _2297_ (.A(_0728_),
    .B(_0729_),
    .C(\reversed_thermometer[164] ),
    .X(_0735_));
 sky130_fd_sc_hd__a221o_1 _2298_ (.A1(\reversed_thermometer[100] ),
    .A2(_0731_),
    .B1(_0732_),
    .B2(\reversed_thermometer[36] ),
    .C1(_0735_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _2299_ (.A(_0728_),
    .B(_0729_),
    .C(\reversed_thermometer[163] ),
    .X(_0736_));
 sky130_fd_sc_hd__a221o_1 _2300_ (.A1(\reversed_thermometer[99] ),
    .A2(_0731_),
    .B1(_0732_),
    .B2(\reversed_thermometer[35] ),
    .C1(_0736_),
    .X(_0256_));
 sky130_fd_sc_hd__buf_1 _2301_ (.A(_0713_),
    .X(_0737_));
 sky130_fd_sc_hd__buf_1 _2302_ (.A(_0715_),
    .X(_0738_));
 sky130_fd_sc_hd__and3_1 _2303_ (.A(_0737_),
    .B(_0738_),
    .C(\reversed_thermometer[162] ),
    .X(_0739_));
 sky130_fd_sc_hd__a221o_1 _2304_ (.A1(\reversed_thermometer[98] ),
    .A2(_0731_),
    .B1(_0732_),
    .B2(\reversed_thermometer[34] ),
    .C1(_0739_),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_2 _2305_ (.A(_0719_),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_2 _2306_ (.A(_0722_),
    .X(_0741_));
 sky130_fd_sc_hd__and3_1 _2307_ (.A(_0737_),
    .B(_0738_),
    .C(\reversed_thermometer[161] ),
    .X(_0742_));
 sky130_fd_sc_hd__a221o_1 _2308_ (.A1(\reversed_thermometer[97] ),
    .A2(_0740_),
    .B1(_0741_),
    .B2(\reversed_thermometer[33] ),
    .C1(_0742_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _2309_ (.A(_0737_),
    .B(_0738_),
    .C(\reversed_thermometer[160] ),
    .X(_0743_));
 sky130_fd_sc_hd__a221o_1 _2310_ (.A1(\reversed_thermometer[96] ),
    .A2(_0740_),
    .B1(_0741_),
    .B2(\reversed_thermometer[32] ),
    .C1(_0743_),
    .X(_0259_));
 sky130_fd_sc_hd__and3_1 _2311_ (.A(_0737_),
    .B(_0738_),
    .C(\reversed_thermometer[159] ),
    .X(_0744_));
 sky130_fd_sc_hd__a221o_1 _2312_ (.A1(\reversed_thermometer[95] ),
    .A2(_0740_),
    .B1(_0741_),
    .B2(\reversed_thermometer[31] ),
    .C1(_0744_),
    .X(_0003_));
 sky130_fd_sc_hd__and3_1 _2313_ (.A(_0737_),
    .B(_0738_),
    .C(\reversed_thermometer[158] ),
    .X(_0745_));
 sky130_fd_sc_hd__a221o_1 _2314_ (.A1(\reversed_thermometer[94] ),
    .A2(_0740_),
    .B1(_0741_),
    .B2(\reversed_thermometer[30] ),
    .C1(_0745_),
    .X(_0004_));
 sky130_fd_sc_hd__buf_1 _2315_ (.A(_0713_),
    .X(_0746_));
 sky130_fd_sc_hd__buf_1 _2316_ (.A(_0715_),
    .X(_0747_));
 sky130_fd_sc_hd__and3_1 _2317_ (.A(_0746_),
    .B(_0747_),
    .C(\reversed_thermometer[157] ),
    .X(_0748_));
 sky130_fd_sc_hd__a221o_1 _2318_ (.A1(\reversed_thermometer[93] ),
    .A2(_0740_),
    .B1(_0741_),
    .B2(\reversed_thermometer[29] ),
    .C1(_0748_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_2 _2319_ (.A(_0719_),
    .X(_0749_));
 sky130_fd_sc_hd__clkbuf_2 _2320_ (.A(_0722_),
    .X(_0750_));
 sky130_fd_sc_hd__and3_1 _2321_ (.A(_0746_),
    .B(_0747_),
    .C(\reversed_thermometer[156] ),
    .X(_0751_));
 sky130_fd_sc_hd__a221o_1 _2322_ (.A1(\reversed_thermometer[92] ),
    .A2(_0749_),
    .B1(_0750_),
    .B2(\reversed_thermometer[28] ),
    .C1(_0751_),
    .X(_0006_));
 sky130_fd_sc_hd__and3_1 _2323_ (.A(_0746_),
    .B(_0747_),
    .C(\reversed_thermometer[155] ),
    .X(_0752_));
 sky130_fd_sc_hd__a221o_1 _2324_ (.A1(\reversed_thermometer[91] ),
    .A2(_0749_),
    .B1(_0750_),
    .B2(\reversed_thermometer[27] ),
    .C1(_0752_),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _2325_ (.A(_0746_),
    .B(_0747_),
    .C(\reversed_thermometer[154] ),
    .X(_0753_));
 sky130_fd_sc_hd__a221o_1 _2326_ (.A1(\reversed_thermometer[90] ),
    .A2(_0749_),
    .B1(_0750_),
    .B2(\reversed_thermometer[26] ),
    .C1(_0753_),
    .X(_0008_));
 sky130_fd_sc_hd__and3_1 _2327_ (.A(_0746_),
    .B(_0747_),
    .C(\reversed_thermometer[153] ),
    .X(_0754_));
 sky130_fd_sc_hd__a221o_1 _2328_ (.A1(\reversed_thermometer[89] ),
    .A2(_0749_),
    .B1(_0750_),
    .B2(\reversed_thermometer[25] ),
    .C1(_0754_),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_2 _2329_ (.A(_0713_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_2 _2330_ (.A(_0715_),
    .X(_0756_));
 sky130_fd_sc_hd__and3_1 _2331_ (.A(_0755_),
    .B(_0756_),
    .C(\reversed_thermometer[152] ),
    .X(_0757_));
 sky130_fd_sc_hd__a221o_1 _2332_ (.A1(\reversed_thermometer[88] ),
    .A2(_0749_),
    .B1(_0750_),
    .B2(\reversed_thermometer[24] ),
    .C1(_0757_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _2333_ (.A(_0719_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_2 _2334_ (.A(_0722_),
    .X(_0759_));
 sky130_fd_sc_hd__and3_1 _2335_ (.A(_0755_),
    .B(_0756_),
    .C(\reversed_thermometer[151] ),
    .X(_0760_));
 sky130_fd_sc_hd__a221o_1 _2336_ (.A1(\reversed_thermometer[87] ),
    .A2(_0758_),
    .B1(_0759_),
    .B2(\reversed_thermometer[23] ),
    .C1(_0760_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _2337_ (.A(_0755_),
    .B(_0756_),
    .C(\reversed_thermometer[150] ),
    .X(_0761_));
 sky130_fd_sc_hd__a221o_1 _2338_ (.A1(\reversed_thermometer[86] ),
    .A2(_0758_),
    .B1(_0759_),
    .B2(\reversed_thermometer[22] ),
    .C1(_0761_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _2339_ (.A(_0755_),
    .B(_0756_),
    .C(\reversed_thermometer[149] ),
    .X(_0762_));
 sky130_fd_sc_hd__a221o_1 _2340_ (.A1(\reversed_thermometer[85] ),
    .A2(_0758_),
    .B1(_0759_),
    .B2(\reversed_thermometer[21] ),
    .C1(_0762_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_1 _2341_ (.A(_0755_),
    .B(_0756_),
    .C(\reversed_thermometer[148] ),
    .X(_0763_));
 sky130_fd_sc_hd__a221o_1 _2342_ (.A1(\reversed_thermometer[84] ),
    .A2(_0758_),
    .B1(_0759_),
    .B2(\reversed_thermometer[20] ),
    .C1(_0763_),
    .X(_0014_));
 sky130_fd_sc_hd__buf_1 _2343_ (.A(\remap_control[0] ),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_4 _2344_ (.A(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__buf_1 _2345_ (.A(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__buf_1 _2346_ (.A(_0670_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_4 _2347_ (.A(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__buf_1 _2348_ (.A(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__and3_1 _2349_ (.A(_0766_),
    .B(_0769_),
    .C(\reversed_thermometer[147] ),
    .X(_0770_));
 sky130_fd_sc_hd__a221o_1 _2350_ (.A1(\reversed_thermometer[83] ),
    .A2(_0758_),
    .B1(_0759_),
    .B2(\reversed_thermometer[19] ),
    .C1(_0770_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _2351_ (.A(_0718_),
    .X(_0771_));
 sky130_fd_sc_hd__clkbuf_2 _2352_ (.A(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _2353_ (.A(_0721_),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_2 _2354_ (.A(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__and3_1 _2355_ (.A(_0766_),
    .B(_0769_),
    .C(\reversed_thermometer[146] ),
    .X(_0775_));
 sky130_fd_sc_hd__a221o_1 _2356_ (.A1(\reversed_thermometer[82] ),
    .A2(_0772_),
    .B1(_0774_),
    .B2(\reversed_thermometer[18] ),
    .C1(_0775_),
    .X(_0016_));
 sky130_fd_sc_hd__and3_1 _2357_ (.A(_0766_),
    .B(_0769_),
    .C(\reversed_thermometer[145] ),
    .X(_0776_));
 sky130_fd_sc_hd__a221o_1 _2358_ (.A1(\reversed_thermometer[81] ),
    .A2(_0772_),
    .B1(_0774_),
    .B2(\reversed_thermometer[17] ),
    .C1(_0776_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _2359_ (.A(_0766_),
    .B(_0769_),
    .C(\reversed_thermometer[144] ),
    .X(_0777_));
 sky130_fd_sc_hd__a221o_1 _2360_ (.A1(\reversed_thermometer[80] ),
    .A2(_0772_),
    .B1(_0774_),
    .B2(\reversed_thermometer[16] ),
    .C1(_0777_),
    .X(_0018_));
 sky130_fd_sc_hd__and3_1 _2361_ (.A(_0766_),
    .B(_0769_),
    .C(\reversed_thermometer[143] ),
    .X(_0778_));
 sky130_fd_sc_hd__a221o_1 _2362_ (.A1(\reversed_thermometer[79] ),
    .A2(_0772_),
    .B1(_0774_),
    .B2(\reversed_thermometer[15] ),
    .C1(_0778_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_1 _2363_ (.A(_0765_),
    .X(_0779_));
 sky130_fd_sc_hd__buf_1 _2364_ (.A(_0768_),
    .X(_0780_));
 sky130_fd_sc_hd__and3_1 _2365_ (.A(_0779_),
    .B(_0780_),
    .C(\reversed_thermometer[142] ),
    .X(_0781_));
 sky130_fd_sc_hd__a221o_1 _2366_ (.A1(\reversed_thermometer[78] ),
    .A2(_0772_),
    .B1(_0774_),
    .B2(\reversed_thermometer[14] ),
    .C1(_0781_),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_2 _2367_ (.A(_0771_),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_2 _2368_ (.A(_0773_),
    .X(_0783_));
 sky130_fd_sc_hd__and3_1 _2369_ (.A(_0779_),
    .B(_0780_),
    .C(\reversed_thermometer[141] ),
    .X(_0784_));
 sky130_fd_sc_hd__a221o_1 _2370_ (.A1(\reversed_thermometer[77] ),
    .A2(_0782_),
    .B1(_0783_),
    .B2(\reversed_thermometer[13] ),
    .C1(_0784_),
    .X(_0021_));
 sky130_fd_sc_hd__and3_1 _2371_ (.A(_0779_),
    .B(_0780_),
    .C(\reversed_thermometer[140] ),
    .X(_0785_));
 sky130_fd_sc_hd__a221o_1 _2372_ (.A1(\reversed_thermometer[76] ),
    .A2(_0782_),
    .B1(_0783_),
    .B2(\reversed_thermometer[12] ),
    .C1(_0785_),
    .X(_0022_));
 sky130_fd_sc_hd__and3_1 _2373_ (.A(_0779_),
    .B(_0780_),
    .C(\reversed_thermometer[139] ),
    .X(_0786_));
 sky130_fd_sc_hd__a221o_1 _2374_ (.A1(\reversed_thermometer[75] ),
    .A2(_0782_),
    .B1(_0783_),
    .B2(\reversed_thermometer[11] ),
    .C1(_0786_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _2375_ (.A(_0779_),
    .B(_0780_),
    .C(\reversed_thermometer[138] ),
    .X(_0787_));
 sky130_fd_sc_hd__a221o_1 _2376_ (.A1(\reversed_thermometer[74] ),
    .A2(_0782_),
    .B1(_0783_),
    .B2(\reversed_thermometer[10] ),
    .C1(_0787_),
    .X(_0024_));
 sky130_fd_sc_hd__buf_1 _2377_ (.A(_0765_),
    .X(_0788_));
 sky130_fd_sc_hd__buf_1 _2378_ (.A(_0768_),
    .X(_0789_));
 sky130_fd_sc_hd__and3_1 _2379_ (.A(_0788_),
    .B(_0789_),
    .C(\reversed_thermometer[137] ),
    .X(_0790_));
 sky130_fd_sc_hd__a221o_1 _2380_ (.A1(\reversed_thermometer[73] ),
    .A2(_0782_),
    .B1(_0783_),
    .B2(\reversed_thermometer[9] ),
    .C1(_0790_),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_2 _2381_ (.A(_0771_),
    .X(_0791_));
 sky130_fd_sc_hd__clkbuf_2 _2382_ (.A(_0773_),
    .X(_0792_));
 sky130_fd_sc_hd__and3_1 _2383_ (.A(_0788_),
    .B(_0789_),
    .C(\reversed_thermometer[136] ),
    .X(_0793_));
 sky130_fd_sc_hd__a221o_1 _2384_ (.A1(\reversed_thermometer[72] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\reversed_thermometer[8] ),
    .C1(_0793_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _2385_ (.A(_0788_),
    .B(_0789_),
    .C(\reversed_thermometer[135] ),
    .X(_0794_));
 sky130_fd_sc_hd__a221o_1 _2386_ (.A1(\reversed_thermometer[71] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\reversed_thermometer[7] ),
    .C1(_0794_),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _2387_ (.A(_0788_),
    .B(_0789_),
    .C(\reversed_thermometer[134] ),
    .X(_0795_));
 sky130_fd_sc_hd__a221o_1 _2388_ (.A1(\reversed_thermometer[70] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\reversed_thermometer[6] ),
    .C1(_0795_),
    .X(_0028_));
 sky130_fd_sc_hd__and3_1 _2389_ (.A(_0788_),
    .B(_0789_),
    .C(\reversed_thermometer[133] ),
    .X(_0796_));
 sky130_fd_sc_hd__a221o_1 _2390_ (.A1(\reversed_thermometer[69] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\reversed_thermometer[5] ),
    .C1(_0796_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_2 _2391_ (.A(_0765_),
    .X(_0797_));
 sky130_fd_sc_hd__clkbuf_2 _2392_ (.A(_0768_),
    .X(_0798_));
 sky130_fd_sc_hd__and3_1 _2393_ (.A(_0797_),
    .B(_0798_),
    .C(\reversed_thermometer[132] ),
    .X(_0799_));
 sky130_fd_sc_hd__a221o_1 _2394_ (.A1(\reversed_thermometer[68] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\reversed_thermometer[4] ),
    .C1(_0799_),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_2 _2395_ (.A(_0771_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_2 _2396_ (.A(_0773_),
    .X(_0801_));
 sky130_fd_sc_hd__and3_1 _2397_ (.A(_0797_),
    .B(_0798_),
    .C(\reversed_thermometer[131] ),
    .X(_0802_));
 sky130_fd_sc_hd__a221o_1 _2398_ (.A1(\reversed_thermometer[67] ),
    .A2(_0800_),
    .B1(_0801_),
    .B2(\reversed_thermometer[3] ),
    .C1(_0802_),
    .X(_0031_));
 sky130_fd_sc_hd__and3_1 _2399_ (.A(_0797_),
    .B(_0798_),
    .C(\reversed_thermometer[130] ),
    .X(_0803_));
 sky130_fd_sc_hd__a221o_1 _2400_ (.A1(\reversed_thermometer[66] ),
    .A2(_0800_),
    .B1(_0801_),
    .B2(\reversed_thermometer[2] ),
    .C1(_0803_),
    .X(_0032_));
 sky130_fd_sc_hd__and3_1 _2401_ (.A(_0797_),
    .B(_0798_),
    .C(\reversed_thermometer[129] ),
    .X(_0804_));
 sky130_fd_sc_hd__a221o_1 _2402_ (.A1(\reversed_thermometer[65] ),
    .A2(_0800_),
    .B1(_0801_),
    .B2(\reversed_thermometer[1] ),
    .C1(_0804_),
    .X(_0033_));
 sky130_fd_sc_hd__and3_1 _2403_ (.A(_0797_),
    .B(_0798_),
    .C(\reversed_thermometer[128] ),
    .X(_0805_));
 sky130_fd_sc_hd__a221o_1 _2404_ (.A1(\reversed_thermometer[64] ),
    .A2(_0800_),
    .B1(_0801_),
    .B2(\reversed_thermometer[0] ),
    .C1(_0805_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_2 _2405_ (.A(_0765_),
    .X(_0806_));
 sky130_fd_sc_hd__clkbuf_2 _2406_ (.A(_0768_),
    .X(_0807_));
 sky130_fd_sc_hd__and3_1 _2407_ (.A(_0806_),
    .B(_0807_),
    .C(\reversed_thermometer[127] ),
    .X(_0808_));
 sky130_fd_sc_hd__a221o_1 _2408_ (.A1(\reversed_thermometer[63] ),
    .A2(_0800_),
    .B1(_0801_),
    .B2(\reversed_thermometer[255] ),
    .C1(_0808_),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_2 _2409_ (.A(_0771_),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_2 _2410_ (.A(_0773_),
    .X(_0810_));
 sky130_fd_sc_hd__and3_1 _2411_ (.A(_0806_),
    .B(_0807_),
    .C(\reversed_thermometer[126] ),
    .X(_0811_));
 sky130_fd_sc_hd__a221o_1 _2412_ (.A1(\reversed_thermometer[62] ),
    .A2(_0809_),
    .B1(_0810_),
    .B2(\reversed_thermometer[254] ),
    .C1(_0811_),
    .X(_0036_));
 sky130_fd_sc_hd__and3_1 _2413_ (.A(_0806_),
    .B(_0807_),
    .C(\reversed_thermometer[125] ),
    .X(_0812_));
 sky130_fd_sc_hd__a221o_1 _2414_ (.A1(\reversed_thermometer[61] ),
    .A2(_0809_),
    .B1(_0810_),
    .B2(\reversed_thermometer[253] ),
    .C1(_0812_),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _2415_ (.A(_0806_),
    .B(_0807_),
    .C(\reversed_thermometer[124] ),
    .X(_0813_));
 sky130_fd_sc_hd__a221o_1 _2416_ (.A1(\reversed_thermometer[60] ),
    .A2(_0809_),
    .B1(_0810_),
    .B2(\reversed_thermometer[252] ),
    .C1(_0813_),
    .X(_0038_));
 sky130_fd_sc_hd__and3_1 _2417_ (.A(_0806_),
    .B(_0807_),
    .C(\reversed_thermometer[123] ),
    .X(_0814_));
 sky130_fd_sc_hd__a221o_1 _2418_ (.A1(\reversed_thermometer[59] ),
    .A2(_0809_),
    .B1(_0810_),
    .B2(\reversed_thermometer[251] ),
    .C1(_0814_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _2419_ (.A(_0764_),
    .X(_0815_));
 sky130_fd_sc_hd__buf_1 _2420_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__buf_2 _2421_ (.A(_0767_),
    .X(_0817_));
 sky130_fd_sc_hd__buf_1 _2422_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__and3_1 _2423_ (.A(_0816_),
    .B(_0818_),
    .C(\reversed_thermometer[122] ),
    .X(_0819_));
 sky130_fd_sc_hd__a221o_1 _2424_ (.A1(\reversed_thermometer[58] ),
    .A2(_0809_),
    .B1(_0810_),
    .B2(\reversed_thermometer[250] ),
    .C1(_0819_),
    .X(_0040_));
 sky130_fd_sc_hd__buf_2 _2425_ (.A(_0718_),
    .X(_0820_));
 sky130_fd_sc_hd__clkbuf_2 _2426_ (.A(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__buf_2 _2427_ (.A(_0721_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_2 _2428_ (.A(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__and3_1 _2429_ (.A(_0816_),
    .B(_0818_),
    .C(\reversed_thermometer[121] ),
    .X(_0824_));
 sky130_fd_sc_hd__a221o_1 _2430_ (.A1(\reversed_thermometer[57] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(\reversed_thermometer[249] ),
    .C1(_0824_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _2431_ (.A(_0816_),
    .B(_0818_),
    .C(\reversed_thermometer[120] ),
    .X(_0825_));
 sky130_fd_sc_hd__a221o_1 _2432_ (.A1(\reversed_thermometer[56] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(\reversed_thermometer[248] ),
    .C1(_0825_),
    .X(_0042_));
 sky130_fd_sc_hd__and3_1 _2433_ (.A(_0816_),
    .B(_0818_),
    .C(\reversed_thermometer[119] ),
    .X(_0826_));
 sky130_fd_sc_hd__a221o_1 _2434_ (.A1(\reversed_thermometer[55] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(\reversed_thermometer[247] ),
    .C1(_0826_),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _2435_ (.A(_0816_),
    .B(_0818_),
    .C(\reversed_thermometer[118] ),
    .X(_0827_));
 sky130_fd_sc_hd__a221o_1 _2436_ (.A1(\reversed_thermometer[54] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(\reversed_thermometer[246] ),
    .C1(_0827_),
    .X(_0044_));
 sky130_fd_sc_hd__buf_1 _2437_ (.A(_0815_),
    .X(_0828_));
 sky130_fd_sc_hd__buf_1 _2438_ (.A(_0817_),
    .X(_0829_));
 sky130_fd_sc_hd__and3_1 _2439_ (.A(_0828_),
    .B(_0829_),
    .C(\reversed_thermometer[117] ),
    .X(_0830_));
 sky130_fd_sc_hd__a221o_1 _2440_ (.A1(\reversed_thermometer[53] ),
    .A2(_0821_),
    .B1(_0823_),
    .B2(\reversed_thermometer[245] ),
    .C1(_0830_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_2 _2441_ (.A(_0820_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_2 _2442_ (.A(_0822_),
    .X(_0832_));
 sky130_fd_sc_hd__and3_1 _2443_ (.A(_0828_),
    .B(_0829_),
    .C(\reversed_thermometer[116] ),
    .X(_0833_));
 sky130_fd_sc_hd__a221o_1 _2444_ (.A1(\reversed_thermometer[52] ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\reversed_thermometer[244] ),
    .C1(_0833_),
    .X(_0046_));
 sky130_fd_sc_hd__and3_1 _2445_ (.A(_0828_),
    .B(_0829_),
    .C(\reversed_thermometer[115] ),
    .X(_0834_));
 sky130_fd_sc_hd__a221o_1 _2446_ (.A1(\reversed_thermometer[51] ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\reversed_thermometer[243] ),
    .C1(_0834_),
    .X(_0047_));
 sky130_fd_sc_hd__and3_1 _2447_ (.A(_0828_),
    .B(_0829_),
    .C(\reversed_thermometer[114] ),
    .X(_0835_));
 sky130_fd_sc_hd__a221o_1 _2448_ (.A1(\reversed_thermometer[50] ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\reversed_thermometer[242] ),
    .C1(_0835_),
    .X(_0048_));
 sky130_fd_sc_hd__and3_1 _2449_ (.A(_0828_),
    .B(_0829_),
    .C(\reversed_thermometer[113] ),
    .X(_0836_));
 sky130_fd_sc_hd__a221o_1 _2450_ (.A1(\reversed_thermometer[49] ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\reversed_thermometer[241] ),
    .C1(_0836_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_1 _2451_ (.A(_0815_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_1 _2452_ (.A(_0817_),
    .X(_0838_));
 sky130_fd_sc_hd__and3_1 _2453_ (.A(_0837_),
    .B(_0838_),
    .C(\reversed_thermometer[112] ),
    .X(_0839_));
 sky130_fd_sc_hd__a221o_1 _2454_ (.A1(\reversed_thermometer[48] ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\reversed_thermometer[240] ),
    .C1(_0839_),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_2 _2455_ (.A(_0820_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_2 _2456_ (.A(_0822_),
    .X(_0841_));
 sky130_fd_sc_hd__and3_1 _2457_ (.A(_0837_),
    .B(_0838_),
    .C(\reversed_thermometer[111] ),
    .X(_0842_));
 sky130_fd_sc_hd__a221o_1 _2458_ (.A1(\reversed_thermometer[47] ),
    .A2(_0840_),
    .B1(_0841_),
    .B2(\reversed_thermometer[239] ),
    .C1(_0842_),
    .X(_0051_));
 sky130_fd_sc_hd__and3_1 _2459_ (.A(_0837_),
    .B(_0838_),
    .C(\reversed_thermometer[110] ),
    .X(_0843_));
 sky130_fd_sc_hd__a221o_1 _2460_ (.A1(\reversed_thermometer[46] ),
    .A2(_0840_),
    .B1(_0841_),
    .B2(\reversed_thermometer[238] ),
    .C1(_0843_),
    .X(_0052_));
 sky130_fd_sc_hd__and3_1 _2461_ (.A(_0837_),
    .B(_0838_),
    .C(\reversed_thermometer[109] ),
    .X(_0844_));
 sky130_fd_sc_hd__a221o_1 _2462_ (.A1(\reversed_thermometer[45] ),
    .A2(_0840_),
    .B1(_0841_),
    .B2(\reversed_thermometer[237] ),
    .C1(_0844_),
    .X(_0053_));
 sky130_fd_sc_hd__and3_1 _2463_ (.A(_0837_),
    .B(_0838_),
    .C(\reversed_thermometer[108] ),
    .X(_0845_));
 sky130_fd_sc_hd__a221o_1 _2464_ (.A1(\reversed_thermometer[44] ),
    .A2(_0840_),
    .B1(_0841_),
    .B2(\reversed_thermometer[236] ),
    .C1(_0845_),
    .X(_0054_));
 sky130_fd_sc_hd__buf_1 _2465_ (.A(_0815_),
    .X(_0846_));
 sky130_fd_sc_hd__buf_1 _2466_ (.A(_0817_),
    .X(_0847_));
 sky130_fd_sc_hd__and3_1 _2467_ (.A(_0846_),
    .B(_0847_),
    .C(\reversed_thermometer[107] ),
    .X(_0848_));
 sky130_fd_sc_hd__a221o_1 _2468_ (.A1(\reversed_thermometer[43] ),
    .A2(_0840_),
    .B1(_0841_),
    .B2(\reversed_thermometer[235] ),
    .C1(_0848_),
    .X(_0055_));
 sky130_fd_sc_hd__clkbuf_2 _2469_ (.A(_0820_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_2 _2470_ (.A(_0822_),
    .X(_0850_));
 sky130_fd_sc_hd__and3_1 _2471_ (.A(_0846_),
    .B(_0847_),
    .C(\reversed_thermometer[106] ),
    .X(_0851_));
 sky130_fd_sc_hd__a221o_1 _2472_ (.A1(\reversed_thermometer[42] ),
    .A2(_0849_),
    .B1(_0850_),
    .B2(\reversed_thermometer[234] ),
    .C1(_0851_),
    .X(_0056_));
 sky130_fd_sc_hd__and3_1 _2473_ (.A(_0846_),
    .B(_0847_),
    .C(\reversed_thermometer[105] ),
    .X(_0852_));
 sky130_fd_sc_hd__a221o_1 _2474_ (.A1(\reversed_thermometer[41] ),
    .A2(_0849_),
    .B1(_0850_),
    .B2(\reversed_thermometer[233] ),
    .C1(_0852_),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _2475_ (.A(_0846_),
    .B(_0847_),
    .C(\reversed_thermometer[104] ),
    .X(_0853_));
 sky130_fd_sc_hd__a221o_1 _2476_ (.A1(\reversed_thermometer[40] ),
    .A2(_0849_),
    .B1(_0850_),
    .B2(\reversed_thermometer[232] ),
    .C1(_0853_),
    .X(_0058_));
 sky130_fd_sc_hd__and3_1 _2477_ (.A(_0846_),
    .B(_0847_),
    .C(\reversed_thermometer[103] ),
    .X(_0854_));
 sky130_fd_sc_hd__a221o_1 _2478_ (.A1(\reversed_thermometer[39] ),
    .A2(_0849_),
    .B1(_0850_),
    .B2(\reversed_thermometer[231] ),
    .C1(_0854_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_1 _2479_ (.A(_0815_),
    .X(_0855_));
 sky130_fd_sc_hd__buf_1 _2480_ (.A(_0817_),
    .X(_0856_));
 sky130_fd_sc_hd__and3_1 _2481_ (.A(_0855_),
    .B(_0856_),
    .C(\reversed_thermometer[102] ),
    .X(_0857_));
 sky130_fd_sc_hd__a221o_1 _2482_ (.A1(\reversed_thermometer[38] ),
    .A2(_0849_),
    .B1(_0850_),
    .B2(\reversed_thermometer[230] ),
    .C1(_0857_),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_2 _2483_ (.A(_0820_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_2 _2484_ (.A(_0822_),
    .X(_0859_));
 sky130_fd_sc_hd__and3_1 _2485_ (.A(_0855_),
    .B(_0856_),
    .C(\reversed_thermometer[101] ),
    .X(_0860_));
 sky130_fd_sc_hd__a221o_1 _2486_ (.A1(\reversed_thermometer[37] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\reversed_thermometer[229] ),
    .C1(_0860_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _2487_ (.A(_0855_),
    .B(_0856_),
    .C(\reversed_thermometer[100] ),
    .X(_0861_));
 sky130_fd_sc_hd__a221o_1 _2488_ (.A1(\reversed_thermometer[36] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\reversed_thermometer[228] ),
    .C1(_0861_),
    .X(_0062_));
 sky130_fd_sc_hd__and3_1 _2489_ (.A(_0855_),
    .B(_0856_),
    .C(\reversed_thermometer[99] ),
    .X(_0862_));
 sky130_fd_sc_hd__a221o_1 _2490_ (.A1(\reversed_thermometer[35] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\reversed_thermometer[227] ),
    .C1(_0862_),
    .X(_0063_));
 sky130_fd_sc_hd__and3_1 _2491_ (.A(_0855_),
    .B(_0856_),
    .C(\reversed_thermometer[98] ),
    .X(_0863_));
 sky130_fd_sc_hd__a221o_1 _2492_ (.A1(\reversed_thermometer[34] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\reversed_thermometer[226] ),
    .C1(_0863_),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_4 _2493_ (.A(_0764_),
    .X(_0864_));
 sky130_fd_sc_hd__buf_1 _2494_ (.A(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_4 _2495_ (.A(_0767_),
    .X(_0866_));
 sky130_fd_sc_hd__buf_1 _2496_ (.A(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__and3_1 _2497_ (.A(_0865_),
    .B(_0867_),
    .C(\reversed_thermometer[97] ),
    .X(_0868_));
 sky130_fd_sc_hd__a221o_1 _2498_ (.A1(\reversed_thermometer[33] ),
    .A2(_0858_),
    .B1(_0859_),
    .B2(\reversed_thermometer[225] ),
    .C1(_0868_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_1 _2499_ (.A(_0674_),
    .X(_0869_));
 sky130_fd_sc_hd__clkbuf_4 _2500_ (.A(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__clkbuf_2 _2501_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__buf_1 _2502_ (.A(_0677_),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_4 _2503_ (.A(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_2 _2504_ (.A(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__and3_1 _2505_ (.A(_0865_),
    .B(_0867_),
    .C(\reversed_thermometer[96] ),
    .X(_0875_));
 sky130_fd_sc_hd__a221o_1 _2506_ (.A1(\reversed_thermometer[32] ),
    .A2(_0871_),
    .B1(_0874_),
    .B2(\reversed_thermometer[224] ),
    .C1(_0875_),
    .X(_0066_));
 sky130_fd_sc_hd__and3_1 _2507_ (.A(_0865_),
    .B(_0867_),
    .C(\reversed_thermometer[95] ),
    .X(_0876_));
 sky130_fd_sc_hd__a221o_1 _2508_ (.A1(\reversed_thermometer[31] ),
    .A2(_0871_),
    .B1(_0874_),
    .B2(\reversed_thermometer[223] ),
    .C1(_0876_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _2509_ (.A(_0865_),
    .B(_0867_),
    .C(\reversed_thermometer[94] ),
    .X(_0877_));
 sky130_fd_sc_hd__a221o_1 _2510_ (.A1(\reversed_thermometer[30] ),
    .A2(_0871_),
    .B1(_0874_),
    .B2(\reversed_thermometer[222] ),
    .C1(_0877_),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _2511_ (.A(_0865_),
    .B(_0867_),
    .C(\reversed_thermometer[93] ),
    .X(_0878_));
 sky130_fd_sc_hd__a221o_1 _2512_ (.A1(\reversed_thermometer[29] ),
    .A2(_0871_),
    .B1(_0874_),
    .B2(\reversed_thermometer[221] ),
    .C1(_0878_),
    .X(_0069_));
 sky130_fd_sc_hd__buf_1 _2513_ (.A(_0864_),
    .X(_0879_));
 sky130_fd_sc_hd__buf_1 _2514_ (.A(_0866_),
    .X(_0880_));
 sky130_fd_sc_hd__and3_1 _2515_ (.A(_0879_),
    .B(_0880_),
    .C(\reversed_thermometer[92] ),
    .X(_0881_));
 sky130_fd_sc_hd__a221o_1 _2516_ (.A1(\reversed_thermometer[28] ),
    .A2(_0871_),
    .B1(_0874_),
    .B2(\reversed_thermometer[220] ),
    .C1(_0881_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_2 _2517_ (.A(_0870_),
    .X(_0882_));
 sky130_fd_sc_hd__clkbuf_2 _2518_ (.A(_0873_),
    .X(_0883_));
 sky130_fd_sc_hd__and3_1 _2519_ (.A(_0879_),
    .B(_0880_),
    .C(\reversed_thermometer[91] ),
    .X(_0884_));
 sky130_fd_sc_hd__a221o_1 _2520_ (.A1(\reversed_thermometer[27] ),
    .A2(_0882_),
    .B1(_0883_),
    .B2(\reversed_thermometer[219] ),
    .C1(_0884_),
    .X(_0071_));
 sky130_fd_sc_hd__and3_1 _2521_ (.A(_0879_),
    .B(_0880_),
    .C(\reversed_thermometer[90] ),
    .X(_0885_));
 sky130_fd_sc_hd__a221o_1 _2522_ (.A1(\reversed_thermometer[26] ),
    .A2(_0882_),
    .B1(_0883_),
    .B2(\reversed_thermometer[218] ),
    .C1(_0885_),
    .X(_0072_));
 sky130_fd_sc_hd__and3_1 _2523_ (.A(_0879_),
    .B(_0880_),
    .C(\reversed_thermometer[89] ),
    .X(_0886_));
 sky130_fd_sc_hd__a221o_1 _2524_ (.A1(\reversed_thermometer[25] ),
    .A2(_0882_),
    .B1(_0883_),
    .B2(\reversed_thermometer[217] ),
    .C1(_0886_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_1 _2525_ (.A(_0879_),
    .B(_0880_),
    .C(\reversed_thermometer[88] ),
    .X(_0887_));
 sky130_fd_sc_hd__a221o_1 _2526_ (.A1(\reversed_thermometer[24] ),
    .A2(_0882_),
    .B1(_0883_),
    .B2(\reversed_thermometer[216] ),
    .C1(_0887_),
    .X(_0074_));
 sky130_fd_sc_hd__buf_1 _2527_ (.A(_0864_),
    .X(_0888_));
 sky130_fd_sc_hd__buf_1 _2528_ (.A(_0866_),
    .X(_0889_));
 sky130_fd_sc_hd__and3_1 _2529_ (.A(_0888_),
    .B(_0889_),
    .C(\reversed_thermometer[87] ),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _2530_ (.A1(\reversed_thermometer[23] ),
    .A2(_0882_),
    .B1(_0883_),
    .B2(\reversed_thermometer[215] ),
    .C1(_0890_),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_2 _2531_ (.A(_0870_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_2 _2532_ (.A(_0873_),
    .X(_0892_));
 sky130_fd_sc_hd__and3_1 _2533_ (.A(_0888_),
    .B(_0889_),
    .C(\reversed_thermometer[86] ),
    .X(_0893_));
 sky130_fd_sc_hd__a221o_1 _2534_ (.A1(\reversed_thermometer[22] ),
    .A2(_0891_),
    .B1(_0892_),
    .B2(\reversed_thermometer[214] ),
    .C1(_0893_),
    .X(_0076_));
 sky130_fd_sc_hd__and3_1 _2535_ (.A(_0888_),
    .B(_0889_),
    .C(\reversed_thermometer[85] ),
    .X(_0894_));
 sky130_fd_sc_hd__a221o_1 _2536_ (.A1(\reversed_thermometer[21] ),
    .A2(_0891_),
    .B1(_0892_),
    .B2(\reversed_thermometer[213] ),
    .C1(_0894_),
    .X(_0077_));
 sky130_fd_sc_hd__and3_1 _2537_ (.A(_0888_),
    .B(_0889_),
    .C(\reversed_thermometer[84] ),
    .X(_0895_));
 sky130_fd_sc_hd__a221o_1 _2538_ (.A1(\reversed_thermometer[20] ),
    .A2(_0891_),
    .B1(_0892_),
    .B2(\reversed_thermometer[212] ),
    .C1(_0895_),
    .X(_0078_));
 sky130_fd_sc_hd__and3_1 _2539_ (.A(_0888_),
    .B(_0889_),
    .C(\reversed_thermometer[83] ),
    .X(_0896_));
 sky130_fd_sc_hd__a221o_1 _2540_ (.A1(\reversed_thermometer[19] ),
    .A2(_0891_),
    .B1(_0892_),
    .B2(\reversed_thermometer[211] ),
    .C1(_0896_),
    .X(_0079_));
 sky130_fd_sc_hd__buf_1 _2541_ (.A(_0864_),
    .X(_0897_));
 sky130_fd_sc_hd__buf_1 _2542_ (.A(_0866_),
    .X(_0898_));
 sky130_fd_sc_hd__and3_1 _2543_ (.A(_0897_),
    .B(_0898_),
    .C(\reversed_thermometer[82] ),
    .X(_0899_));
 sky130_fd_sc_hd__a221o_1 _2544_ (.A1(\reversed_thermometer[18] ),
    .A2(_0891_),
    .B1(_0892_),
    .B2(\reversed_thermometer[210] ),
    .C1(_0899_),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_2 _2545_ (.A(_0870_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_2 _2546_ (.A(_0873_),
    .X(_0901_));
 sky130_fd_sc_hd__and3_1 _2547_ (.A(_0897_),
    .B(_0898_),
    .C(\reversed_thermometer[81] ),
    .X(_0902_));
 sky130_fd_sc_hd__a221o_1 _2548_ (.A1(\reversed_thermometer[17] ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\reversed_thermometer[209] ),
    .C1(_0902_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _2549_ (.A(_0897_),
    .B(_0898_),
    .C(\reversed_thermometer[80] ),
    .X(_0903_));
 sky130_fd_sc_hd__a221o_1 _2550_ (.A1(\reversed_thermometer[16] ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\reversed_thermometer[208] ),
    .C1(_0903_),
    .X(_0082_));
 sky130_fd_sc_hd__and3_1 _2551_ (.A(_0897_),
    .B(_0898_),
    .C(\reversed_thermometer[79] ),
    .X(_0904_));
 sky130_fd_sc_hd__a221o_1 _2552_ (.A1(\reversed_thermometer[15] ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\reversed_thermometer[207] ),
    .C1(_0904_),
    .X(_0083_));
 sky130_fd_sc_hd__and3_1 _2553_ (.A(_0897_),
    .B(_0898_),
    .C(\reversed_thermometer[78] ),
    .X(_0905_));
 sky130_fd_sc_hd__a221o_1 _2554_ (.A1(\reversed_thermometer[14] ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\reversed_thermometer[206] ),
    .C1(_0905_),
    .X(_0084_));
 sky130_fd_sc_hd__buf_1 _2555_ (.A(_0864_),
    .X(_0906_));
 sky130_fd_sc_hd__buf_1 _2556_ (.A(_0866_),
    .X(_0907_));
 sky130_fd_sc_hd__and3_1 _2557_ (.A(_0906_),
    .B(_0907_),
    .C(\reversed_thermometer[77] ),
    .X(_0908_));
 sky130_fd_sc_hd__a221o_1 _2558_ (.A1(\reversed_thermometer[13] ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\reversed_thermometer[205] ),
    .C1(_0908_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_2 _2559_ (.A(_0870_),
    .X(_0909_));
 sky130_fd_sc_hd__clkbuf_2 _2560_ (.A(_0873_),
    .X(_0910_));
 sky130_fd_sc_hd__and3_1 _2561_ (.A(_0906_),
    .B(_0907_),
    .C(\reversed_thermometer[76] ),
    .X(_0911_));
 sky130_fd_sc_hd__a221o_1 _2562_ (.A1(\reversed_thermometer[12] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(\reversed_thermometer[204] ),
    .C1(_0911_),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _2563_ (.A(_0906_),
    .B(_0907_),
    .C(\reversed_thermometer[75] ),
    .X(_0912_));
 sky130_fd_sc_hd__a221o_1 _2564_ (.A1(\reversed_thermometer[11] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(\reversed_thermometer[203] ),
    .C1(_0912_),
    .X(_0087_));
 sky130_fd_sc_hd__and3_1 _2565_ (.A(_0906_),
    .B(_0907_),
    .C(\reversed_thermometer[74] ),
    .X(_0913_));
 sky130_fd_sc_hd__a221o_1 _2566_ (.A1(\reversed_thermometer[10] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(\reversed_thermometer[202] ),
    .C1(_0913_),
    .X(_0088_));
 sky130_fd_sc_hd__and3_1 _2567_ (.A(_0906_),
    .B(_0907_),
    .C(\reversed_thermometer[73] ),
    .X(_0914_));
 sky130_fd_sc_hd__a221o_1 _2568_ (.A1(\reversed_thermometer[9] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(\reversed_thermometer[201] ),
    .C1(_0914_),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_4 _2569_ (.A(_0764_),
    .X(_0915_));
 sky130_fd_sc_hd__buf_1 _2570_ (.A(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__clkbuf_4 _2571_ (.A(_0767_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_2 _2572_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__and3_1 _2573_ (.A(_0916_),
    .B(_0918_),
    .C(\reversed_thermometer[72] ),
    .X(_0919_));
 sky130_fd_sc_hd__a221o_1 _2574_ (.A1(\reversed_thermometer[8] ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(\reversed_thermometer[200] ),
    .C1(_0919_),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_2 _2575_ (.A(_0869_),
    .X(_0920_));
 sky130_fd_sc_hd__buf_2 _2576_ (.A(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_2 _2577_ (.A(_0872_),
    .X(_0922_));
 sky130_fd_sc_hd__buf_2 _2578_ (.A(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__and3_1 _2579_ (.A(_0916_),
    .B(_0918_),
    .C(\reversed_thermometer[71] ),
    .X(_0924_));
 sky130_fd_sc_hd__a221o_1 _2580_ (.A1(\reversed_thermometer[7] ),
    .A2(_0921_),
    .B1(_0923_),
    .B2(\reversed_thermometer[199] ),
    .C1(_0924_),
    .X(_0091_));
 sky130_fd_sc_hd__and3_1 _2581_ (.A(_0916_),
    .B(_0918_),
    .C(\reversed_thermometer[70] ),
    .X(_0925_));
 sky130_fd_sc_hd__a221o_1 _2582_ (.A1(\reversed_thermometer[6] ),
    .A2(_0921_),
    .B1(_0923_),
    .B2(\reversed_thermometer[198] ),
    .C1(_0925_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _2583_ (.A(_0916_),
    .B(_0918_),
    .C(\reversed_thermometer[69] ),
    .X(_0926_));
 sky130_fd_sc_hd__a221o_1 _2584_ (.A1(\reversed_thermometer[5] ),
    .A2(_0921_),
    .B1(_0923_),
    .B2(\reversed_thermometer[197] ),
    .C1(_0926_),
    .X(_0093_));
 sky130_fd_sc_hd__and3_1 _2585_ (.A(_0916_),
    .B(_0918_),
    .C(\reversed_thermometer[68] ),
    .X(_0927_));
 sky130_fd_sc_hd__a221o_1 _2586_ (.A1(\reversed_thermometer[4] ),
    .A2(_0921_),
    .B1(_0923_),
    .B2(\reversed_thermometer[196] ),
    .C1(_0927_),
    .X(_0094_));
 sky130_fd_sc_hd__buf_1 _2587_ (.A(_0915_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_2 _2588_ (.A(_0917_),
    .X(_0929_));
 sky130_fd_sc_hd__and3_1 _2589_ (.A(_0928_),
    .B(_0929_),
    .C(\reversed_thermometer[67] ),
    .X(_0930_));
 sky130_fd_sc_hd__a221o_1 _2590_ (.A1(\reversed_thermometer[3] ),
    .A2(_0921_),
    .B1(_0923_),
    .B2(\reversed_thermometer[195] ),
    .C1(_0930_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_2 _2591_ (.A(_0920_),
    .X(_0931_));
 sky130_fd_sc_hd__buf_2 _2592_ (.A(_0922_),
    .X(_0932_));
 sky130_fd_sc_hd__and3_1 _2593_ (.A(_0928_),
    .B(_0929_),
    .C(\reversed_thermometer[66] ),
    .X(_0933_));
 sky130_fd_sc_hd__a221o_1 _2594_ (.A1(\reversed_thermometer[2] ),
    .A2(_0931_),
    .B1(_0932_),
    .B2(\reversed_thermometer[194] ),
    .C1(_0933_),
    .X(_0096_));
 sky130_fd_sc_hd__and3_1 _2595_ (.A(_0928_),
    .B(_0929_),
    .C(\reversed_thermometer[65] ),
    .X(_0934_));
 sky130_fd_sc_hd__a221o_1 _2596_ (.A1(\reversed_thermometer[1] ),
    .A2(_0931_),
    .B1(_0932_),
    .B2(\reversed_thermometer[193] ),
    .C1(_0934_),
    .X(_0097_));
 sky130_fd_sc_hd__and3_1 _2597_ (.A(_0928_),
    .B(_0929_),
    .C(\reversed_thermometer[64] ),
    .X(_0935_));
 sky130_fd_sc_hd__a221o_1 _2598_ (.A1(\reversed_thermometer[0] ),
    .A2(_0931_),
    .B1(_0932_),
    .B2(\reversed_thermometer[192] ),
    .C1(_0935_),
    .X(_0098_));
 sky130_fd_sc_hd__and3_1 _2599_ (.A(_0928_),
    .B(_0929_),
    .C(\reversed_thermometer[63] ),
    .X(_0936_));
 sky130_fd_sc_hd__a221o_1 _2600_ (.A1(\reversed_thermometer[255] ),
    .A2(_0931_),
    .B1(_0932_),
    .B2(\reversed_thermometer[191] ),
    .C1(_0936_),
    .X(_0099_));
 sky130_fd_sc_hd__buf_1 _2601_ (.A(_0915_),
    .X(_0937_));
 sky130_fd_sc_hd__buf_1 _2602_ (.A(_0917_),
    .X(_0938_));
 sky130_fd_sc_hd__and3_1 _2603_ (.A(_0937_),
    .B(_0938_),
    .C(\reversed_thermometer[62] ),
    .X(_0939_));
 sky130_fd_sc_hd__a221o_1 _2604_ (.A1(\reversed_thermometer[254] ),
    .A2(_0931_),
    .B1(_0932_),
    .B2(\reversed_thermometer[190] ),
    .C1(_0939_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_2 _2605_ (.A(_0920_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_2 _2606_ (.A(_0922_),
    .X(_0941_));
 sky130_fd_sc_hd__and3_1 _2607_ (.A(_0937_),
    .B(_0938_),
    .C(\reversed_thermometer[61] ),
    .X(_0942_));
 sky130_fd_sc_hd__a221o_1 _2608_ (.A1(\reversed_thermometer[253] ),
    .A2(_0940_),
    .B1(_0941_),
    .B2(\reversed_thermometer[189] ),
    .C1(_0942_),
    .X(_0101_));
 sky130_fd_sc_hd__and3_1 _2609_ (.A(_0937_),
    .B(_0938_),
    .C(\reversed_thermometer[60] ),
    .X(_0943_));
 sky130_fd_sc_hd__a221o_1 _2610_ (.A1(\reversed_thermometer[252] ),
    .A2(_0940_),
    .B1(_0941_),
    .B2(\reversed_thermometer[188] ),
    .C1(_0943_),
    .X(_0102_));
 sky130_fd_sc_hd__and3_1 _2611_ (.A(_0937_),
    .B(_0938_),
    .C(\reversed_thermometer[59] ),
    .X(_0944_));
 sky130_fd_sc_hd__a221o_1 _2612_ (.A1(\reversed_thermometer[251] ),
    .A2(_0940_),
    .B1(_0941_),
    .B2(\reversed_thermometer[187] ),
    .C1(_0944_),
    .X(_0103_));
 sky130_fd_sc_hd__and3_1 _2613_ (.A(_0937_),
    .B(_0938_),
    .C(\reversed_thermometer[58] ),
    .X(_0945_));
 sky130_fd_sc_hd__a221o_1 _2614_ (.A1(\reversed_thermometer[250] ),
    .A2(_0940_),
    .B1(_0941_),
    .B2(\reversed_thermometer[186] ),
    .C1(_0945_),
    .X(_0104_));
 sky130_fd_sc_hd__buf_1 _2615_ (.A(_0915_),
    .X(_0946_));
 sky130_fd_sc_hd__buf_1 _2616_ (.A(_0917_),
    .X(_0947_));
 sky130_fd_sc_hd__and3_1 _2617_ (.A(_0946_),
    .B(_0947_),
    .C(\reversed_thermometer[57] ),
    .X(_0948_));
 sky130_fd_sc_hd__a221o_1 _2618_ (.A1(\reversed_thermometer[249] ),
    .A2(_0940_),
    .B1(_0941_),
    .B2(\reversed_thermometer[185] ),
    .C1(_0948_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_2 _2619_ (.A(_0920_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_2 _2620_ (.A(_0922_),
    .X(_0950_));
 sky130_fd_sc_hd__and3_1 _2621_ (.A(_0946_),
    .B(_0947_),
    .C(\reversed_thermometer[56] ),
    .X(_0951_));
 sky130_fd_sc_hd__a221o_1 _2622_ (.A1(\reversed_thermometer[248] ),
    .A2(_0949_),
    .B1(_0950_),
    .B2(\reversed_thermometer[184] ),
    .C1(_0951_),
    .X(_0106_));
 sky130_fd_sc_hd__and3_1 _2623_ (.A(_0946_),
    .B(_0947_),
    .C(\reversed_thermometer[55] ),
    .X(_0952_));
 sky130_fd_sc_hd__a221o_1 _2624_ (.A1(\reversed_thermometer[247] ),
    .A2(_0949_),
    .B1(_0950_),
    .B2(\reversed_thermometer[183] ),
    .C1(_0952_),
    .X(_0107_));
 sky130_fd_sc_hd__and3_1 _2625_ (.A(_0946_),
    .B(_0947_),
    .C(\reversed_thermometer[54] ),
    .X(_0953_));
 sky130_fd_sc_hd__a221o_1 _2626_ (.A1(\reversed_thermometer[246] ),
    .A2(_0949_),
    .B1(_0950_),
    .B2(\reversed_thermometer[182] ),
    .C1(_0953_),
    .X(_0108_));
 sky130_fd_sc_hd__and3_1 _2627_ (.A(_0946_),
    .B(_0947_),
    .C(\reversed_thermometer[53] ),
    .X(_0954_));
 sky130_fd_sc_hd__a221o_1 _2628_ (.A1(\reversed_thermometer[245] ),
    .A2(_0949_),
    .B1(_0950_),
    .B2(\reversed_thermometer[181] ),
    .C1(_0954_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_1 _2629_ (.A(_0915_),
    .X(_0955_));
 sky130_fd_sc_hd__buf_1 _2630_ (.A(_0917_),
    .X(_0956_));
 sky130_fd_sc_hd__and3_1 _2631_ (.A(_0955_),
    .B(_0956_),
    .C(\reversed_thermometer[52] ),
    .X(_0957_));
 sky130_fd_sc_hd__a221o_1 _2632_ (.A1(\reversed_thermometer[244] ),
    .A2(_0949_),
    .B1(_0950_),
    .B2(\reversed_thermometer[180] ),
    .C1(_0957_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_2 _2633_ (.A(_0920_),
    .X(_0958_));
 sky130_fd_sc_hd__clkbuf_2 _2634_ (.A(_0922_),
    .X(_0959_));
 sky130_fd_sc_hd__and3_1 _2635_ (.A(_0955_),
    .B(_0956_),
    .C(\reversed_thermometer[51] ),
    .X(_0960_));
 sky130_fd_sc_hd__a221o_1 _2636_ (.A1(\reversed_thermometer[243] ),
    .A2(_0958_),
    .B1(_0959_),
    .B2(\reversed_thermometer[179] ),
    .C1(_0960_),
    .X(_0111_));
 sky130_fd_sc_hd__and3_1 _2637_ (.A(_0955_),
    .B(_0956_),
    .C(\reversed_thermometer[50] ),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _2638_ (.A1(\reversed_thermometer[242] ),
    .A2(_0958_),
    .B1(_0959_),
    .B2(\reversed_thermometer[178] ),
    .C1(_0961_),
    .X(_0112_));
 sky130_fd_sc_hd__and3_1 _2639_ (.A(_0955_),
    .B(_0956_),
    .C(\reversed_thermometer[49] ),
    .X(_0962_));
 sky130_fd_sc_hd__a221o_1 _2640_ (.A1(\reversed_thermometer[241] ),
    .A2(_0958_),
    .B1(_0959_),
    .B2(\reversed_thermometer[177] ),
    .C1(_0962_),
    .X(_0113_));
 sky130_fd_sc_hd__and3_1 _2641_ (.A(_0955_),
    .B(_0956_),
    .C(\reversed_thermometer[48] ),
    .X(_0963_));
 sky130_fd_sc_hd__a221o_1 _2642_ (.A1(\reversed_thermometer[240] ),
    .A2(_0958_),
    .B1(_0959_),
    .B2(\reversed_thermometer[176] ),
    .C1(_0963_),
    .X(_0114_));
 sky130_fd_sc_hd__buf_2 _2643_ (.A(_0764_),
    .X(_0964_));
 sky130_fd_sc_hd__buf_1 _2644_ (.A(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__buf_2 _2645_ (.A(_0767_),
    .X(_0966_));
 sky130_fd_sc_hd__buf_1 _2646_ (.A(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__and3_1 _2647_ (.A(_0965_),
    .B(_0967_),
    .C(\reversed_thermometer[47] ),
    .X(_0968_));
 sky130_fd_sc_hd__a221o_1 _2648_ (.A1(\reversed_thermometer[239] ),
    .A2(_0958_),
    .B1(_0959_),
    .B2(\reversed_thermometer[175] ),
    .C1(_0968_),
    .X(_0115_));
 sky130_fd_sc_hd__buf_2 _2649_ (.A(_0869_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_2 _2650_ (.A(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__buf_2 _2651_ (.A(_0872_),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_2 _2652_ (.A(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__and3_1 _2653_ (.A(_0965_),
    .B(_0967_),
    .C(\reversed_thermometer[46] ),
    .X(_0973_));
 sky130_fd_sc_hd__a221o_1 _2654_ (.A1(\reversed_thermometer[238] ),
    .A2(_0970_),
    .B1(_0972_),
    .B2(\reversed_thermometer[174] ),
    .C1(_0973_),
    .X(_0116_));
 sky130_fd_sc_hd__and3_1 _2655_ (.A(_0965_),
    .B(_0967_),
    .C(\reversed_thermometer[45] ),
    .X(_0974_));
 sky130_fd_sc_hd__a221o_1 _2656_ (.A1(\reversed_thermometer[237] ),
    .A2(_0970_),
    .B1(_0972_),
    .B2(\reversed_thermometer[173] ),
    .C1(_0974_),
    .X(_0117_));
 sky130_fd_sc_hd__and3_1 _2657_ (.A(_0965_),
    .B(_0967_),
    .C(\reversed_thermometer[44] ),
    .X(_0975_));
 sky130_fd_sc_hd__a221o_1 _2658_ (.A1(\reversed_thermometer[236] ),
    .A2(_0970_),
    .B1(_0972_),
    .B2(\reversed_thermometer[172] ),
    .C1(_0975_),
    .X(_0118_));
 sky130_fd_sc_hd__and3_1 _2659_ (.A(_0965_),
    .B(_0967_),
    .C(\reversed_thermometer[43] ),
    .X(_0976_));
 sky130_fd_sc_hd__a221o_1 _2660_ (.A1(\reversed_thermometer[235] ),
    .A2(_0970_),
    .B1(_0972_),
    .B2(\reversed_thermometer[171] ),
    .C1(_0976_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_1 _2661_ (.A(_0964_),
    .X(_0977_));
 sky130_fd_sc_hd__buf_1 _2662_ (.A(_0966_),
    .X(_0978_));
 sky130_fd_sc_hd__and3_1 _2663_ (.A(_0977_),
    .B(_0978_),
    .C(\reversed_thermometer[42] ),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _2664_ (.A1(\reversed_thermometer[234] ),
    .A2(_0970_),
    .B1(_0972_),
    .B2(\reversed_thermometer[170] ),
    .C1(_0979_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_2 _2665_ (.A(_0969_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_2 _2666_ (.A(_0971_),
    .X(_0981_));
 sky130_fd_sc_hd__and3_1 _2667_ (.A(_0977_),
    .B(_0978_),
    .C(\reversed_thermometer[41] ),
    .X(_0982_));
 sky130_fd_sc_hd__a221o_1 _2668_ (.A1(\reversed_thermometer[233] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\reversed_thermometer[169] ),
    .C1(_0982_),
    .X(_0121_));
 sky130_fd_sc_hd__and3_1 _2669_ (.A(_0977_),
    .B(_0978_),
    .C(\reversed_thermometer[40] ),
    .X(_0983_));
 sky130_fd_sc_hd__a221o_1 _2670_ (.A1(\reversed_thermometer[232] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\reversed_thermometer[168] ),
    .C1(_0983_),
    .X(_0122_));
 sky130_fd_sc_hd__and3_1 _2671_ (.A(_0977_),
    .B(_0978_),
    .C(\reversed_thermometer[39] ),
    .X(_0984_));
 sky130_fd_sc_hd__a221o_1 _2672_ (.A1(\reversed_thermometer[231] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\reversed_thermometer[167] ),
    .C1(_0984_),
    .X(_0123_));
 sky130_fd_sc_hd__and3_1 _2673_ (.A(_0977_),
    .B(_0978_),
    .C(\reversed_thermometer[38] ),
    .X(_0985_));
 sky130_fd_sc_hd__a221o_1 _2674_ (.A1(\reversed_thermometer[230] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\reversed_thermometer[166] ),
    .C1(_0985_),
    .X(_0124_));
 sky130_fd_sc_hd__buf_1 _2675_ (.A(_0964_),
    .X(_0986_));
 sky130_fd_sc_hd__buf_1 _2676_ (.A(_0966_),
    .X(_0987_));
 sky130_fd_sc_hd__and3_1 _2677_ (.A(_0986_),
    .B(_0987_),
    .C(\reversed_thermometer[37] ),
    .X(_0988_));
 sky130_fd_sc_hd__a221o_1 _2678_ (.A1(\reversed_thermometer[229] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\reversed_thermometer[165] ),
    .C1(_0988_),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_2 _2679_ (.A(_0969_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_2 _2680_ (.A(_0971_),
    .X(_0990_));
 sky130_fd_sc_hd__and3_1 _2681_ (.A(_0986_),
    .B(_0987_),
    .C(\reversed_thermometer[36] ),
    .X(_0991_));
 sky130_fd_sc_hd__a221o_1 _2682_ (.A1(\reversed_thermometer[228] ),
    .A2(_0989_),
    .B1(_0990_),
    .B2(\reversed_thermometer[164] ),
    .C1(_0991_),
    .X(_0126_));
 sky130_fd_sc_hd__and3_1 _2683_ (.A(_0986_),
    .B(_0987_),
    .C(\reversed_thermometer[35] ),
    .X(_0992_));
 sky130_fd_sc_hd__a221o_1 _2684_ (.A1(\reversed_thermometer[227] ),
    .A2(_0989_),
    .B1(_0990_),
    .B2(\reversed_thermometer[163] ),
    .C1(_0992_),
    .X(_0127_));
 sky130_fd_sc_hd__and3_1 _2685_ (.A(_0986_),
    .B(_0987_),
    .C(\reversed_thermometer[34] ),
    .X(_0993_));
 sky130_fd_sc_hd__a221o_1 _2686_ (.A1(\reversed_thermometer[226] ),
    .A2(_0989_),
    .B1(_0990_),
    .B2(\reversed_thermometer[162] ),
    .C1(_0993_),
    .X(_0128_));
 sky130_fd_sc_hd__and3_1 _2687_ (.A(_0986_),
    .B(_0987_),
    .C(\reversed_thermometer[33] ),
    .X(_0994_));
 sky130_fd_sc_hd__a221o_1 _2688_ (.A1(\reversed_thermometer[225] ),
    .A2(_0989_),
    .B1(_0990_),
    .B2(\reversed_thermometer[161] ),
    .C1(_0994_),
    .X(_0129_));
 sky130_fd_sc_hd__buf_1 _2689_ (.A(_0964_),
    .X(_0995_));
 sky130_fd_sc_hd__buf_1 _2690_ (.A(_0966_),
    .X(_0996_));
 sky130_fd_sc_hd__and3_1 _2691_ (.A(_0995_),
    .B(_0996_),
    .C(\reversed_thermometer[32] ),
    .X(_0997_));
 sky130_fd_sc_hd__a221o_1 _2692_ (.A1(\reversed_thermometer[224] ),
    .A2(_0989_),
    .B1(_0990_),
    .B2(\reversed_thermometer[160] ),
    .C1(_0997_),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_2 _2693_ (.A(_0969_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_2 _2694_ (.A(_0971_),
    .X(_0999_));
 sky130_fd_sc_hd__and3_1 _2695_ (.A(_0995_),
    .B(_0996_),
    .C(\reversed_thermometer[31] ),
    .X(_1000_));
 sky130_fd_sc_hd__a221o_1 _2696_ (.A1(\reversed_thermometer[223] ),
    .A2(_0998_),
    .B1(_0999_),
    .B2(\reversed_thermometer[159] ),
    .C1(_1000_),
    .X(_0131_));
 sky130_fd_sc_hd__and3_1 _2697_ (.A(_0995_),
    .B(_0996_),
    .C(\reversed_thermometer[30] ),
    .X(_1001_));
 sky130_fd_sc_hd__a221o_1 _2698_ (.A1(\reversed_thermometer[222] ),
    .A2(_0998_),
    .B1(_0999_),
    .B2(\reversed_thermometer[158] ),
    .C1(_1001_),
    .X(_0132_));
 sky130_fd_sc_hd__and3_1 _2699_ (.A(_0995_),
    .B(_0996_),
    .C(\reversed_thermometer[29] ),
    .X(_1002_));
 sky130_fd_sc_hd__a221o_1 _2700_ (.A1(\reversed_thermometer[221] ),
    .A2(_0998_),
    .B1(_0999_),
    .B2(\reversed_thermometer[157] ),
    .C1(_1002_),
    .X(_0133_));
 sky130_fd_sc_hd__and3_1 _2701_ (.A(_0995_),
    .B(_0996_),
    .C(\reversed_thermometer[28] ),
    .X(_1003_));
 sky130_fd_sc_hd__a221o_1 _2702_ (.A1(\reversed_thermometer[220] ),
    .A2(_0998_),
    .B1(_0999_),
    .B2(\reversed_thermometer[156] ),
    .C1(_1003_),
    .X(_0134_));
 sky130_fd_sc_hd__buf_1 _2703_ (.A(_0964_),
    .X(_1004_));
 sky130_fd_sc_hd__buf_1 _2704_ (.A(_0966_),
    .X(_1005_));
 sky130_fd_sc_hd__and3_1 _2705_ (.A(_1004_),
    .B(_1005_),
    .C(\reversed_thermometer[27] ),
    .X(_1006_));
 sky130_fd_sc_hd__a221o_1 _2706_ (.A1(\reversed_thermometer[219] ),
    .A2(_0998_),
    .B1(_0999_),
    .B2(\reversed_thermometer[155] ),
    .C1(_1006_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_2 _2707_ (.A(_0969_),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_2 _2708_ (.A(_0971_),
    .X(_1008_));
 sky130_fd_sc_hd__and3_1 _2709_ (.A(_1004_),
    .B(_1005_),
    .C(\reversed_thermometer[26] ),
    .X(_1009_));
 sky130_fd_sc_hd__a221o_1 _2710_ (.A1(\reversed_thermometer[218] ),
    .A2(_1007_),
    .B1(_1008_),
    .B2(\reversed_thermometer[154] ),
    .C1(_1009_),
    .X(_0136_));
 sky130_fd_sc_hd__and3_1 _2711_ (.A(_1004_),
    .B(_1005_),
    .C(\reversed_thermometer[25] ),
    .X(_1010_));
 sky130_fd_sc_hd__a221o_1 _2712_ (.A1(\reversed_thermometer[217] ),
    .A2(_1007_),
    .B1(_1008_),
    .B2(\reversed_thermometer[153] ),
    .C1(_1010_),
    .X(_0137_));
 sky130_fd_sc_hd__and3_1 _2713_ (.A(_1004_),
    .B(_1005_),
    .C(\reversed_thermometer[24] ),
    .X(_1011_));
 sky130_fd_sc_hd__a221o_1 _2714_ (.A1(\reversed_thermometer[216] ),
    .A2(_1007_),
    .B1(_1008_),
    .B2(\reversed_thermometer[152] ),
    .C1(_1011_),
    .X(_0138_));
 sky130_fd_sc_hd__and3_1 _2715_ (.A(_1004_),
    .B(_1005_),
    .C(\reversed_thermometer[23] ),
    .X(_1012_));
 sky130_fd_sc_hd__a221o_1 _2716_ (.A1(\reversed_thermometer[215] ),
    .A2(_1007_),
    .B1(_1008_),
    .B2(\reversed_thermometer[151] ),
    .C1(_1012_),
    .X(_0139_));
 sky130_fd_sc_hd__buf_2 _2717_ (.A(_0667_),
    .X(_1013_));
 sky130_fd_sc_hd__buf_1 _2718_ (.A(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__buf_2 _2719_ (.A(_0670_),
    .X(_1015_));
 sky130_fd_sc_hd__buf_1 _2720_ (.A(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__and3_1 _2721_ (.A(_1014_),
    .B(_1016_),
    .C(\reversed_thermometer[22] ),
    .X(_1017_));
 sky130_fd_sc_hd__a221o_1 _2722_ (.A1(\reversed_thermometer[214] ),
    .A2(_1007_),
    .B1(_1008_),
    .B2(\reversed_thermometer[150] ),
    .C1(_1017_),
    .X(_0140_));
 sky130_fd_sc_hd__buf_2 _2723_ (.A(_0869_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_2 _2724_ (.A(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__buf_2 _2725_ (.A(_0872_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_2 _2726_ (.A(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__and3_1 _2727_ (.A(_1014_),
    .B(_1016_),
    .C(\reversed_thermometer[21] ),
    .X(_1022_));
 sky130_fd_sc_hd__a221o_1 _2728_ (.A1(\reversed_thermometer[213] ),
    .A2(_1019_),
    .B1(_1021_),
    .B2(\reversed_thermometer[149] ),
    .C1(_1022_),
    .X(_0141_));
 sky130_fd_sc_hd__and3_1 _2729_ (.A(_1014_),
    .B(_1016_),
    .C(\reversed_thermometer[20] ),
    .X(_1023_));
 sky130_fd_sc_hd__a221o_1 _2730_ (.A1(\reversed_thermometer[212] ),
    .A2(_1019_),
    .B1(_1021_),
    .B2(\reversed_thermometer[148] ),
    .C1(_1023_),
    .X(_0142_));
 sky130_fd_sc_hd__and3_1 _2731_ (.A(_1014_),
    .B(_1016_),
    .C(\reversed_thermometer[19] ),
    .X(_1024_));
 sky130_fd_sc_hd__a221o_1 _2732_ (.A1(\reversed_thermometer[211] ),
    .A2(_1019_),
    .B1(_1021_),
    .B2(\reversed_thermometer[147] ),
    .C1(_1024_),
    .X(_0143_));
 sky130_fd_sc_hd__and3_1 _2733_ (.A(_1014_),
    .B(_1016_),
    .C(\reversed_thermometer[18] ),
    .X(_1025_));
 sky130_fd_sc_hd__a221o_1 _2734_ (.A1(\reversed_thermometer[210] ),
    .A2(_1019_),
    .B1(_1021_),
    .B2(\reversed_thermometer[146] ),
    .C1(_1025_),
    .X(_0144_));
 sky130_fd_sc_hd__buf_1 _2735_ (.A(_1013_),
    .X(_1026_));
 sky130_fd_sc_hd__buf_1 _2736_ (.A(_1015_),
    .X(_1027_));
 sky130_fd_sc_hd__and3_1 _2737_ (.A(_1026_),
    .B(_1027_),
    .C(\reversed_thermometer[17] ),
    .X(_1028_));
 sky130_fd_sc_hd__a221o_1 _2738_ (.A1(\reversed_thermometer[209] ),
    .A2(_1019_),
    .B1(_1021_),
    .B2(\reversed_thermometer[145] ),
    .C1(_1028_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_2 _2739_ (.A(_1018_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_2 _2740_ (.A(_1020_),
    .X(_1030_));
 sky130_fd_sc_hd__and3_1 _2741_ (.A(_1026_),
    .B(_1027_),
    .C(\reversed_thermometer[16] ),
    .X(_1031_));
 sky130_fd_sc_hd__a221o_1 _2742_ (.A1(\reversed_thermometer[208] ),
    .A2(_1029_),
    .B1(_1030_),
    .B2(\reversed_thermometer[144] ),
    .C1(_1031_),
    .X(_0146_));
 sky130_fd_sc_hd__and3_1 _2743_ (.A(_1026_),
    .B(_1027_),
    .C(\reversed_thermometer[15] ),
    .X(_1032_));
 sky130_fd_sc_hd__a221o_1 _2744_ (.A1(\reversed_thermometer[207] ),
    .A2(_1029_),
    .B1(_1030_),
    .B2(\reversed_thermometer[143] ),
    .C1(_1032_),
    .X(_0147_));
 sky130_fd_sc_hd__and3_1 _2745_ (.A(_1026_),
    .B(_1027_),
    .C(\reversed_thermometer[14] ),
    .X(_1033_));
 sky130_fd_sc_hd__a221o_1 _2746_ (.A1(\reversed_thermometer[206] ),
    .A2(_1029_),
    .B1(_1030_),
    .B2(\reversed_thermometer[142] ),
    .C1(_1033_),
    .X(_0148_));
 sky130_fd_sc_hd__and3_1 _2747_ (.A(_1026_),
    .B(_1027_),
    .C(\reversed_thermometer[13] ),
    .X(_1034_));
 sky130_fd_sc_hd__a221o_1 _2748_ (.A1(\reversed_thermometer[205] ),
    .A2(_1029_),
    .B1(_1030_),
    .B2(\reversed_thermometer[141] ),
    .C1(_1034_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_1 _2749_ (.A(_1013_),
    .X(_1035_));
 sky130_fd_sc_hd__buf_1 _2750_ (.A(_1015_),
    .X(_1036_));
 sky130_fd_sc_hd__and3_1 _2751_ (.A(_1035_),
    .B(_1036_),
    .C(\reversed_thermometer[12] ),
    .X(_1037_));
 sky130_fd_sc_hd__a221o_1 _2752_ (.A1(\reversed_thermometer[204] ),
    .A2(_1029_),
    .B1(_1030_),
    .B2(\reversed_thermometer[140] ),
    .C1(_1037_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_2 _2753_ (.A(_1018_),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_2 _2754_ (.A(_1020_),
    .X(_1039_));
 sky130_fd_sc_hd__and3_1 _2755_ (.A(_1035_),
    .B(_1036_),
    .C(\reversed_thermometer[11] ),
    .X(_1040_));
 sky130_fd_sc_hd__a221o_1 _2756_ (.A1(\reversed_thermometer[203] ),
    .A2(_1038_),
    .B1(_1039_),
    .B2(\reversed_thermometer[139] ),
    .C1(_1040_),
    .X(_0151_));
 sky130_fd_sc_hd__and3_1 _2757_ (.A(_1035_),
    .B(_1036_),
    .C(\reversed_thermometer[10] ),
    .X(_1041_));
 sky130_fd_sc_hd__a221o_1 _2758_ (.A1(\reversed_thermometer[202] ),
    .A2(_1038_),
    .B1(_1039_),
    .B2(\reversed_thermometer[138] ),
    .C1(_1041_),
    .X(_0152_));
 sky130_fd_sc_hd__and3_1 _2759_ (.A(_1035_),
    .B(_1036_),
    .C(\reversed_thermometer[9] ),
    .X(_1042_));
 sky130_fd_sc_hd__a221o_1 _2760_ (.A1(\reversed_thermometer[201] ),
    .A2(_1038_),
    .B1(_1039_),
    .B2(\reversed_thermometer[137] ),
    .C1(_1042_),
    .X(_0153_));
 sky130_fd_sc_hd__and3_1 _2761_ (.A(_1035_),
    .B(_1036_),
    .C(\reversed_thermometer[8] ),
    .X(_1043_));
 sky130_fd_sc_hd__a221o_1 _2762_ (.A1(\reversed_thermometer[200] ),
    .A2(_1038_),
    .B1(_1039_),
    .B2(\reversed_thermometer[136] ),
    .C1(_1043_),
    .X(_0154_));
 sky130_fd_sc_hd__buf_1 _2763_ (.A(_1013_),
    .X(_1044_));
 sky130_fd_sc_hd__buf_1 _2764_ (.A(_1015_),
    .X(_1045_));
 sky130_fd_sc_hd__and3_1 _2765_ (.A(_1044_),
    .B(_1045_),
    .C(\reversed_thermometer[7] ),
    .X(_1046_));
 sky130_fd_sc_hd__a221o_1 _2766_ (.A1(\reversed_thermometer[199] ),
    .A2(_1038_),
    .B1(_1039_),
    .B2(\reversed_thermometer[135] ),
    .C1(_1046_),
    .X(_0155_));
 sky130_fd_sc_hd__buf_2 _2767_ (.A(_1018_),
    .X(_1047_));
 sky130_fd_sc_hd__buf_2 _2768_ (.A(_1020_),
    .X(_1048_));
 sky130_fd_sc_hd__and3_1 _2769_ (.A(_1044_),
    .B(_1045_),
    .C(\reversed_thermometer[6] ),
    .X(_1049_));
 sky130_fd_sc_hd__a221o_1 _2770_ (.A1(\reversed_thermometer[198] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(\reversed_thermometer[134] ),
    .C1(_1049_),
    .X(_0156_));
 sky130_fd_sc_hd__and3_1 _2771_ (.A(_1044_),
    .B(_1045_),
    .C(\reversed_thermometer[5] ),
    .X(_1050_));
 sky130_fd_sc_hd__a221o_1 _2772_ (.A1(\reversed_thermometer[197] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(\reversed_thermometer[133] ),
    .C1(_1050_),
    .X(_0157_));
 sky130_fd_sc_hd__and3_1 _2773_ (.A(_1044_),
    .B(_1045_),
    .C(\reversed_thermometer[4] ),
    .X(_1051_));
 sky130_fd_sc_hd__a221o_1 _2774_ (.A1(\reversed_thermometer[196] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(\reversed_thermometer[132] ),
    .C1(_1051_),
    .X(_0158_));
 sky130_fd_sc_hd__and3_1 _2775_ (.A(_1044_),
    .B(_1045_),
    .C(\reversed_thermometer[3] ),
    .X(_1052_));
 sky130_fd_sc_hd__a221o_1 _2776_ (.A1(\reversed_thermometer[195] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(\reversed_thermometer[131] ),
    .C1(_1052_),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_2 _2777_ (.A(_1013_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_2 _2778_ (.A(_1015_),
    .X(_1054_));
 sky130_fd_sc_hd__and3_1 _2779_ (.A(_1053_),
    .B(_1054_),
    .C(\reversed_thermometer[2] ),
    .X(_1055_));
 sky130_fd_sc_hd__a221o_1 _2780_ (.A1(\reversed_thermometer[194] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(\reversed_thermometer[130] ),
    .C1(_1055_),
    .X(_0160_));
 sky130_fd_sc_hd__buf_2 _2781_ (.A(_1018_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_2 _2782_ (.A(_1020_),
    .X(_1057_));
 sky130_fd_sc_hd__and3_1 _2783_ (.A(_1053_),
    .B(_1054_),
    .C(\reversed_thermometer[1] ),
    .X(_1058_));
 sky130_fd_sc_hd__a221o_1 _2784_ (.A1(\reversed_thermometer[193] ),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\reversed_thermometer[129] ),
    .C1(_1058_),
    .X(_0161_));
 sky130_fd_sc_hd__and3_1 _2785_ (.A(_1053_),
    .B(_1054_),
    .C(\reversed_thermometer[0] ),
    .X(_1059_));
 sky130_fd_sc_hd__a221o_1 _2786_ (.A1(\reversed_thermometer[192] ),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\reversed_thermometer[128] ),
    .C1(_1059_),
    .X(_0162_));
 sky130_fd_sc_hd__and3_1 _2787_ (.A(_1053_),
    .B(_1054_),
    .C(\reversed_thermometer[255] ),
    .X(_1060_));
 sky130_fd_sc_hd__a221o_1 _2788_ (.A1(\reversed_thermometer[191] ),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\reversed_thermometer[127] ),
    .C1(_1060_),
    .X(_0163_));
 sky130_fd_sc_hd__and3_1 _2789_ (.A(_1053_),
    .B(_1054_),
    .C(\reversed_thermometer[254] ),
    .X(_1061_));
 sky130_fd_sc_hd__a221o_1 _2790_ (.A1(\reversed_thermometer[190] ),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\reversed_thermometer[126] ),
    .C1(_1061_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_4 _2791_ (.A(_0667_),
    .X(_1062_));
 sky130_fd_sc_hd__buf_1 _2792_ (.A(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_4 _2793_ (.A(_0670_),
    .X(_1064_));
 sky130_fd_sc_hd__buf_1 _2794_ (.A(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__and3_1 _2795_ (.A(_1063_),
    .B(_1065_),
    .C(\reversed_thermometer[253] ),
    .X(_1066_));
 sky130_fd_sc_hd__a221o_1 _2796_ (.A1(\reversed_thermometer[189] ),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\reversed_thermometer[125] ),
    .C1(_1066_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _2797_ (.A(_0869_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_2 _2798_ (.A(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__buf_2 _2799_ (.A(_0872_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_2 _2800_ (.A(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__and3_1 _2801_ (.A(_1063_),
    .B(_1065_),
    .C(\reversed_thermometer[252] ),
    .X(_1071_));
 sky130_fd_sc_hd__a221o_1 _2802_ (.A1(\reversed_thermometer[188] ),
    .A2(_1068_),
    .B1(_1070_),
    .B2(\reversed_thermometer[124] ),
    .C1(_1071_),
    .X(_0166_));
 sky130_fd_sc_hd__and3_1 _2803_ (.A(_1063_),
    .B(_1065_),
    .C(\reversed_thermometer[251] ),
    .X(_1072_));
 sky130_fd_sc_hd__a221o_1 _2804_ (.A1(\reversed_thermometer[187] ),
    .A2(_1068_),
    .B1(_1070_),
    .B2(\reversed_thermometer[123] ),
    .C1(_1072_),
    .X(_0167_));
 sky130_fd_sc_hd__and3_1 _2805_ (.A(_1063_),
    .B(_1065_),
    .C(\reversed_thermometer[250] ),
    .X(_1073_));
 sky130_fd_sc_hd__a221o_1 _2806_ (.A1(\reversed_thermometer[186] ),
    .A2(_1068_),
    .B1(_1070_),
    .B2(\reversed_thermometer[122] ),
    .C1(_1073_),
    .X(_0168_));
 sky130_fd_sc_hd__and3_1 _2807_ (.A(_1063_),
    .B(_1065_),
    .C(\reversed_thermometer[249] ),
    .X(_1074_));
 sky130_fd_sc_hd__a221o_1 _2808_ (.A1(\reversed_thermometer[185] ),
    .A2(_1068_),
    .B1(_1070_),
    .B2(\reversed_thermometer[121] ),
    .C1(_1074_),
    .X(_0169_));
 sky130_fd_sc_hd__buf_1 _2809_ (.A(_1062_),
    .X(_1075_));
 sky130_fd_sc_hd__buf_1 _2810_ (.A(_1064_),
    .X(_1076_));
 sky130_fd_sc_hd__and3_1 _2811_ (.A(_1075_),
    .B(_1076_),
    .C(\reversed_thermometer[248] ),
    .X(_1077_));
 sky130_fd_sc_hd__a221o_1 _2812_ (.A1(\reversed_thermometer[184] ),
    .A2(_1068_),
    .B1(_1070_),
    .B2(\reversed_thermometer[120] ),
    .C1(_1077_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_2 _2813_ (.A(_1067_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_2 _2814_ (.A(_1069_),
    .X(_1079_));
 sky130_fd_sc_hd__and3_1 _2815_ (.A(_1075_),
    .B(_1076_),
    .C(\reversed_thermometer[247] ),
    .X(_1080_));
 sky130_fd_sc_hd__a221o_1 _2816_ (.A1(\reversed_thermometer[183] ),
    .A2(_1078_),
    .B1(_1079_),
    .B2(\reversed_thermometer[119] ),
    .C1(_1080_),
    .X(_0171_));
 sky130_fd_sc_hd__and3_1 _2817_ (.A(_1075_),
    .B(_1076_),
    .C(\reversed_thermometer[246] ),
    .X(_1081_));
 sky130_fd_sc_hd__a221o_1 _2818_ (.A1(\reversed_thermometer[182] ),
    .A2(_1078_),
    .B1(_1079_),
    .B2(\reversed_thermometer[118] ),
    .C1(_1081_),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _2819_ (.A(_1075_),
    .B(_1076_),
    .C(\reversed_thermometer[245] ),
    .X(_1082_));
 sky130_fd_sc_hd__a221o_1 _2820_ (.A1(\reversed_thermometer[181] ),
    .A2(_1078_),
    .B1(_1079_),
    .B2(\reversed_thermometer[117] ),
    .C1(_1082_),
    .X(_0173_));
 sky130_fd_sc_hd__and3_1 _2821_ (.A(_1075_),
    .B(_1076_),
    .C(\reversed_thermometer[244] ),
    .X(_1083_));
 sky130_fd_sc_hd__a221o_1 _2822_ (.A1(\reversed_thermometer[180] ),
    .A2(_1078_),
    .B1(_1079_),
    .B2(\reversed_thermometer[116] ),
    .C1(_1083_),
    .X(_0174_));
 sky130_fd_sc_hd__buf_1 _2823_ (.A(_1062_),
    .X(_1084_));
 sky130_fd_sc_hd__buf_1 _2824_ (.A(_1064_),
    .X(_1085_));
 sky130_fd_sc_hd__and3_1 _2825_ (.A(_1084_),
    .B(_1085_),
    .C(\reversed_thermometer[243] ),
    .X(_1086_));
 sky130_fd_sc_hd__a221o_1 _2826_ (.A1(\reversed_thermometer[179] ),
    .A2(_1078_),
    .B1(_1079_),
    .B2(\reversed_thermometer[115] ),
    .C1(_1086_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_2 _2827_ (.A(_1067_),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_2 _2828_ (.A(_1069_),
    .X(_1088_));
 sky130_fd_sc_hd__and3_1 _2829_ (.A(_1084_),
    .B(_1085_),
    .C(\reversed_thermometer[242] ),
    .X(_1089_));
 sky130_fd_sc_hd__a221o_1 _2830_ (.A1(\reversed_thermometer[178] ),
    .A2(_1087_),
    .B1(_1088_),
    .B2(\reversed_thermometer[114] ),
    .C1(_1089_),
    .X(_0176_));
 sky130_fd_sc_hd__and3_1 _2831_ (.A(_1084_),
    .B(_1085_),
    .C(\reversed_thermometer[241] ),
    .X(_1090_));
 sky130_fd_sc_hd__a221o_1 _2832_ (.A1(\reversed_thermometer[177] ),
    .A2(_1087_),
    .B1(_1088_),
    .B2(\reversed_thermometer[113] ),
    .C1(_1090_),
    .X(_0177_));
 sky130_fd_sc_hd__and3_1 _2833_ (.A(_1084_),
    .B(_1085_),
    .C(\reversed_thermometer[240] ),
    .X(_1091_));
 sky130_fd_sc_hd__a221o_1 _2834_ (.A1(\reversed_thermometer[176] ),
    .A2(_1087_),
    .B1(_1088_),
    .B2(\reversed_thermometer[112] ),
    .C1(_1091_),
    .X(_0178_));
 sky130_fd_sc_hd__and3_1 _2835_ (.A(_1084_),
    .B(_1085_),
    .C(\reversed_thermometer[239] ),
    .X(_1092_));
 sky130_fd_sc_hd__a221o_1 _2836_ (.A1(\reversed_thermometer[175] ),
    .A2(_1087_),
    .B1(_1088_),
    .B2(\reversed_thermometer[111] ),
    .C1(_1092_),
    .X(_0179_));
 sky130_fd_sc_hd__buf_1 _2837_ (.A(_1062_),
    .X(_1093_));
 sky130_fd_sc_hd__buf_1 _2838_ (.A(_1064_),
    .X(_1094_));
 sky130_fd_sc_hd__and3_1 _2839_ (.A(_1093_),
    .B(_1094_),
    .C(\reversed_thermometer[238] ),
    .X(_1095_));
 sky130_fd_sc_hd__a221o_1 _2840_ (.A1(\reversed_thermometer[174] ),
    .A2(_1087_),
    .B1(_1088_),
    .B2(\reversed_thermometer[110] ),
    .C1(_1095_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_2 _2841_ (.A(_1067_),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_2 _2842_ (.A(_1069_),
    .X(_1097_));
 sky130_fd_sc_hd__and3_1 _2843_ (.A(_1093_),
    .B(_1094_),
    .C(\reversed_thermometer[237] ),
    .X(_1098_));
 sky130_fd_sc_hd__a221o_1 _2844_ (.A1(\reversed_thermometer[173] ),
    .A2(_1096_),
    .B1(_1097_),
    .B2(\reversed_thermometer[109] ),
    .C1(_1098_),
    .X(_0181_));
 sky130_fd_sc_hd__and3_1 _2845_ (.A(_1093_),
    .B(_1094_),
    .C(\reversed_thermometer[236] ),
    .X(_1099_));
 sky130_fd_sc_hd__a221o_1 _2846_ (.A1(\reversed_thermometer[172] ),
    .A2(_1096_),
    .B1(_1097_),
    .B2(\reversed_thermometer[108] ),
    .C1(_1099_),
    .X(_0182_));
 sky130_fd_sc_hd__and3_1 _2847_ (.A(_1093_),
    .B(_1094_),
    .C(\reversed_thermometer[235] ),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _2848_ (.A1(\reversed_thermometer[171] ),
    .A2(_1096_),
    .B1(_1097_),
    .B2(\reversed_thermometer[107] ),
    .C1(_1100_),
    .X(_0183_));
 sky130_fd_sc_hd__and3_1 _2849_ (.A(_1093_),
    .B(_1094_),
    .C(\reversed_thermometer[234] ),
    .X(_1101_));
 sky130_fd_sc_hd__a221o_1 _2850_ (.A1(\reversed_thermometer[170] ),
    .A2(_1096_),
    .B1(_1097_),
    .B2(\reversed_thermometer[106] ),
    .C1(_1101_),
    .X(_0184_));
 sky130_fd_sc_hd__buf_1 _2851_ (.A(_1062_),
    .X(_1102_));
 sky130_fd_sc_hd__buf_1 _2852_ (.A(_1064_),
    .X(_1103_));
 sky130_fd_sc_hd__and3_1 _2853_ (.A(_1102_),
    .B(_1103_),
    .C(\reversed_thermometer[233] ),
    .X(_1104_));
 sky130_fd_sc_hd__a221o_1 _2854_ (.A1(\reversed_thermometer[169] ),
    .A2(_1096_),
    .B1(_1097_),
    .B2(\reversed_thermometer[105] ),
    .C1(_1104_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_2 _2855_ (.A(_1067_),
    .X(_1105_));
 sky130_fd_sc_hd__clkbuf_2 _2856_ (.A(_1069_),
    .X(_1106_));
 sky130_fd_sc_hd__and3_1 _2857_ (.A(_1102_),
    .B(_1103_),
    .C(\reversed_thermometer[232] ),
    .X(_1107_));
 sky130_fd_sc_hd__a221o_1 _2858_ (.A1(\reversed_thermometer[168] ),
    .A2(_1105_),
    .B1(_1106_),
    .B2(\reversed_thermometer[104] ),
    .C1(_1107_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _2859_ (.A(_1102_),
    .B(_1103_),
    .C(\reversed_thermometer[231] ),
    .X(_1108_));
 sky130_fd_sc_hd__a221o_1 _2860_ (.A1(\reversed_thermometer[167] ),
    .A2(_1105_),
    .B1(_1106_),
    .B2(\reversed_thermometer[103] ),
    .C1(_1108_),
    .X(_0187_));
 sky130_fd_sc_hd__and3_1 _2861_ (.A(_1102_),
    .B(_1103_),
    .C(\reversed_thermometer[230] ),
    .X(_1109_));
 sky130_fd_sc_hd__a221o_1 _2862_ (.A1(\reversed_thermometer[166] ),
    .A2(_1105_),
    .B1(_1106_),
    .B2(\reversed_thermometer[102] ),
    .C1(_1109_),
    .X(_0188_));
 sky130_fd_sc_hd__and3_1 _2863_ (.A(_1102_),
    .B(_1103_),
    .C(\reversed_thermometer[229] ),
    .X(_1110_));
 sky130_fd_sc_hd__a221o_1 _2864_ (.A1(\reversed_thermometer[165] ),
    .A2(_1105_),
    .B1(_1106_),
    .B2(\reversed_thermometer[101] ),
    .C1(_1110_),
    .X(_0189_));
 sky130_fd_sc_hd__buf_2 _2865_ (.A(_0667_),
    .X(_1111_));
 sky130_fd_sc_hd__buf_1 _2866_ (.A(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__buf_2 _2867_ (.A(_0670_),
    .X(_1113_));
 sky130_fd_sc_hd__buf_1 _2868_ (.A(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__and3_1 _2869_ (.A(_1112_),
    .B(_1114_),
    .C(\reversed_thermometer[228] ),
    .X(_1115_));
 sky130_fd_sc_hd__a221o_1 _2870_ (.A1(\reversed_thermometer[164] ),
    .A2(_1105_),
    .B1(_1106_),
    .B2(\reversed_thermometer[100] ),
    .C1(_1115_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_4 _2871_ (.A(_0674_),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_2 _2872_ (.A(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_4 _2873_ (.A(_0677_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_2 _2874_ (.A(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__and3_1 _2875_ (.A(_1112_),
    .B(_1114_),
    .C(\reversed_thermometer[227] ),
    .X(_1120_));
 sky130_fd_sc_hd__a221o_1 _2876_ (.A1(\reversed_thermometer[163] ),
    .A2(_1117_),
    .B1(_1119_),
    .B2(\reversed_thermometer[99] ),
    .C1(_1120_),
    .X(_0191_));
 sky130_fd_sc_hd__and3_1 _2877_ (.A(_1112_),
    .B(_1114_),
    .C(\reversed_thermometer[226] ),
    .X(_1121_));
 sky130_fd_sc_hd__a221o_1 _2878_ (.A1(\reversed_thermometer[162] ),
    .A2(_1117_),
    .B1(_1119_),
    .B2(\reversed_thermometer[98] ),
    .C1(_1121_),
    .X(_0192_));
 sky130_fd_sc_hd__and3_1 _2879_ (.A(_1112_),
    .B(_1114_),
    .C(\reversed_thermometer[225] ),
    .X(_1122_));
 sky130_fd_sc_hd__a221o_1 _2880_ (.A1(\reversed_thermometer[161] ),
    .A2(_1117_),
    .B1(_1119_),
    .B2(\reversed_thermometer[97] ),
    .C1(_1122_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_1 _2881_ (.A(_1112_),
    .B(_1114_),
    .C(\reversed_thermometer[224] ),
    .X(_1123_));
 sky130_fd_sc_hd__a221o_1 _2882_ (.A1(\reversed_thermometer[160] ),
    .A2(_1117_),
    .B1(_1119_),
    .B2(\reversed_thermometer[96] ),
    .C1(_1123_),
    .X(_0194_));
 sky130_fd_sc_hd__buf_1 _2883_ (.A(_1111_),
    .X(_1124_));
 sky130_fd_sc_hd__buf_1 _2884_ (.A(_1113_),
    .X(_1125_));
 sky130_fd_sc_hd__and3_1 _2885_ (.A(_1124_),
    .B(_1125_),
    .C(\reversed_thermometer[223] ),
    .X(_1126_));
 sky130_fd_sc_hd__a221o_1 _2886_ (.A1(\reversed_thermometer[159] ),
    .A2(_1117_),
    .B1(_1119_),
    .B2(\reversed_thermometer[95] ),
    .C1(_1126_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_2 _2887_ (.A(_1116_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_2 _2888_ (.A(_1118_),
    .X(_1128_));
 sky130_fd_sc_hd__and3_1 _2889_ (.A(_1124_),
    .B(_1125_),
    .C(\reversed_thermometer[222] ),
    .X(_1129_));
 sky130_fd_sc_hd__a221o_1 _2890_ (.A1(\reversed_thermometer[158] ),
    .A2(_1127_),
    .B1(_1128_),
    .B2(\reversed_thermometer[94] ),
    .C1(_1129_),
    .X(_0196_));
 sky130_fd_sc_hd__and3_1 _2891_ (.A(_1124_),
    .B(_1125_),
    .C(\reversed_thermometer[221] ),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_1 _2892_ (.A1(\reversed_thermometer[157] ),
    .A2(_1127_),
    .B1(_1128_),
    .B2(\reversed_thermometer[93] ),
    .C1(_1130_),
    .X(_0197_));
 sky130_fd_sc_hd__and3_1 _2893_ (.A(_1124_),
    .B(_1125_),
    .C(\reversed_thermometer[220] ),
    .X(_1131_));
 sky130_fd_sc_hd__a221o_1 _2894_ (.A1(\reversed_thermometer[156] ),
    .A2(_1127_),
    .B1(_1128_),
    .B2(\reversed_thermometer[92] ),
    .C1(_1131_),
    .X(_0198_));
 sky130_fd_sc_hd__and3_1 _2895_ (.A(_1124_),
    .B(_1125_),
    .C(\reversed_thermometer[219] ),
    .X(_1132_));
 sky130_fd_sc_hd__a221o_1 _2896_ (.A1(\reversed_thermometer[155] ),
    .A2(_1127_),
    .B1(_1128_),
    .B2(\reversed_thermometer[91] ),
    .C1(_1132_),
    .X(_0199_));
 sky130_fd_sc_hd__buf_1 _2897_ (.A(_1111_),
    .X(_1133_));
 sky130_fd_sc_hd__buf_1 _2898_ (.A(_1113_),
    .X(_1134_));
 sky130_fd_sc_hd__and3_1 _2899_ (.A(_1133_),
    .B(_1134_),
    .C(\reversed_thermometer[218] ),
    .X(_1135_));
 sky130_fd_sc_hd__a221o_1 _2900_ (.A1(\reversed_thermometer[154] ),
    .A2(_1127_),
    .B1(_1128_),
    .B2(\reversed_thermometer[90] ),
    .C1(_1135_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_2 _2901_ (.A(_1116_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_2 _2902_ (.A(_1118_),
    .X(_1137_));
 sky130_fd_sc_hd__and3_1 _2903_ (.A(_1133_),
    .B(_1134_),
    .C(\reversed_thermometer[217] ),
    .X(_1138_));
 sky130_fd_sc_hd__a221o_1 _2904_ (.A1(\reversed_thermometer[153] ),
    .A2(_1136_),
    .B1(_1137_),
    .B2(\reversed_thermometer[89] ),
    .C1(_1138_),
    .X(_0201_));
 sky130_fd_sc_hd__and3_1 _2905_ (.A(_1133_),
    .B(_1134_),
    .C(\reversed_thermometer[216] ),
    .X(_1139_));
 sky130_fd_sc_hd__a221o_1 _2906_ (.A1(\reversed_thermometer[152] ),
    .A2(_1136_),
    .B1(_1137_),
    .B2(\reversed_thermometer[88] ),
    .C1(_1139_),
    .X(_0202_));
 sky130_fd_sc_hd__and3_1 _2907_ (.A(_1133_),
    .B(_1134_),
    .C(\reversed_thermometer[215] ),
    .X(_1140_));
 sky130_fd_sc_hd__a221o_1 _2908_ (.A1(\reversed_thermometer[151] ),
    .A2(_1136_),
    .B1(_1137_),
    .B2(\reversed_thermometer[87] ),
    .C1(_1140_),
    .X(_0203_));
 sky130_fd_sc_hd__and3_1 _2909_ (.A(_1133_),
    .B(_1134_),
    .C(\reversed_thermometer[214] ),
    .X(_1141_));
 sky130_fd_sc_hd__a221o_1 _2910_ (.A1(\reversed_thermometer[150] ),
    .A2(_1136_),
    .B1(_1137_),
    .B2(\reversed_thermometer[86] ),
    .C1(_1141_),
    .X(_0204_));
 sky130_fd_sc_hd__buf_1 _2911_ (.A(_1111_),
    .X(_1142_));
 sky130_fd_sc_hd__buf_1 _2912_ (.A(_1113_),
    .X(_1143_));
 sky130_fd_sc_hd__and3_1 _2913_ (.A(_1142_),
    .B(_1143_),
    .C(\reversed_thermometer[213] ),
    .X(_1144_));
 sky130_fd_sc_hd__a221o_1 _2914_ (.A1(\reversed_thermometer[149] ),
    .A2(_1136_),
    .B1(_1137_),
    .B2(\reversed_thermometer[85] ),
    .C1(_1144_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_2 _2915_ (.A(_1116_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_2 _2916_ (.A(_1118_),
    .X(_1146_));
 sky130_fd_sc_hd__and3_1 _2917_ (.A(_1142_),
    .B(_1143_),
    .C(\reversed_thermometer[212] ),
    .X(_1147_));
 sky130_fd_sc_hd__a221o_1 _2918_ (.A1(\reversed_thermometer[148] ),
    .A2(_1145_),
    .B1(_1146_),
    .B2(\reversed_thermometer[84] ),
    .C1(_1147_),
    .X(_0206_));
 sky130_fd_sc_hd__and3_1 _2919_ (.A(_1142_),
    .B(_1143_),
    .C(\reversed_thermometer[211] ),
    .X(_1148_));
 sky130_fd_sc_hd__a221o_1 _2920_ (.A1(\reversed_thermometer[147] ),
    .A2(_1145_),
    .B1(_1146_),
    .B2(\reversed_thermometer[83] ),
    .C1(_1148_),
    .X(_0207_));
 sky130_fd_sc_hd__and3_1 _2921_ (.A(_1142_),
    .B(_1143_),
    .C(\reversed_thermometer[210] ),
    .X(_1149_));
 sky130_fd_sc_hd__a221o_1 _2922_ (.A1(\reversed_thermometer[146] ),
    .A2(_1145_),
    .B1(_1146_),
    .B2(\reversed_thermometer[82] ),
    .C1(_1149_),
    .X(_0208_));
 sky130_fd_sc_hd__and3_1 _2923_ (.A(_1142_),
    .B(_1143_),
    .C(\reversed_thermometer[209] ),
    .X(_1150_));
 sky130_fd_sc_hd__a221o_1 _2924_ (.A1(\reversed_thermometer[145] ),
    .A2(_1145_),
    .B1(_1146_),
    .B2(\reversed_thermometer[81] ),
    .C1(_1150_),
    .X(_0209_));
 sky130_fd_sc_hd__buf_1 _2925_ (.A(_1111_),
    .X(_1151_));
 sky130_fd_sc_hd__buf_1 _2926_ (.A(_1113_),
    .X(_1152_));
 sky130_fd_sc_hd__and3_1 _2927_ (.A(_1151_),
    .B(_1152_),
    .C(\reversed_thermometer[208] ),
    .X(_1153_));
 sky130_fd_sc_hd__a221o_1 _2928_ (.A1(\reversed_thermometer[144] ),
    .A2(_1145_),
    .B1(_1146_),
    .B2(\reversed_thermometer[80] ),
    .C1(_1153_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_2 _2929_ (.A(_1116_),
    .X(_1154_));
 sky130_fd_sc_hd__clkbuf_2 _2930_ (.A(_1118_),
    .X(_1155_));
 sky130_fd_sc_hd__and3_1 _2931_ (.A(_1151_),
    .B(_1152_),
    .C(\reversed_thermometer[207] ),
    .X(_1156_));
 sky130_fd_sc_hd__a221o_1 _2932_ (.A1(\reversed_thermometer[143] ),
    .A2(_1154_),
    .B1(_1155_),
    .B2(\reversed_thermometer[79] ),
    .C1(_1156_),
    .X(_0211_));
 sky130_fd_sc_hd__and3_1 _2933_ (.A(_1151_),
    .B(_1152_),
    .C(\reversed_thermometer[206] ),
    .X(_1157_));
 sky130_fd_sc_hd__a221o_1 _2934_ (.A1(\reversed_thermometer[142] ),
    .A2(_1154_),
    .B1(_1155_),
    .B2(\reversed_thermometer[78] ),
    .C1(_1157_),
    .X(_0212_));
 sky130_fd_sc_hd__and3_1 _2935_ (.A(_1151_),
    .B(_1152_),
    .C(\reversed_thermometer[205] ),
    .X(_1158_));
 sky130_fd_sc_hd__a221o_1 _2936_ (.A1(\reversed_thermometer[141] ),
    .A2(_1154_),
    .B1(_1155_),
    .B2(\reversed_thermometer[77] ),
    .C1(_1158_),
    .X(_0213_));
 sky130_fd_sc_hd__and3_1 _2937_ (.A(_1151_),
    .B(_1152_),
    .C(\reversed_thermometer[204] ),
    .X(_1159_));
 sky130_fd_sc_hd__a221o_1 _2938_ (.A1(\reversed_thermometer[140] ),
    .A2(_1154_),
    .B1(_1155_),
    .B2(\reversed_thermometer[76] ),
    .C1(_1159_),
    .X(_0214_));
 sky130_fd_sc_hd__buf_1 _2939_ (.A(_0668_),
    .X(_1160_));
 sky130_fd_sc_hd__buf_1 _2940_ (.A(_0671_),
    .X(_1161_));
 sky130_fd_sc_hd__and3_1 _2941_ (.A(_1160_),
    .B(_1161_),
    .C(\reversed_thermometer[203] ),
    .X(_1162_));
 sky130_fd_sc_hd__a221o_1 _2942_ (.A1(\reversed_thermometer[139] ),
    .A2(_1154_),
    .B1(_1155_),
    .B2(\reversed_thermometer[75] ),
    .C1(_1162_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_2 _2943_ (.A(_0718_),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_2 _2944_ (.A(_0721_),
    .X(_1164_));
 sky130_fd_sc_hd__and3_1 _2945_ (.A(_1160_),
    .B(_1161_),
    .C(\reversed_thermometer[202] ),
    .X(_1165_));
 sky130_fd_sc_hd__a221o_1 _2946_ (.A1(\reversed_thermometer[138] ),
    .A2(_1163_),
    .B1(_1164_),
    .B2(\reversed_thermometer[74] ),
    .C1(_1165_),
    .X(_0216_));
 sky130_fd_sc_hd__and3_1 _2947_ (.A(_1160_),
    .B(_1161_),
    .C(\reversed_thermometer[201] ),
    .X(_1166_));
 sky130_fd_sc_hd__a221o_1 _2948_ (.A1(\reversed_thermometer[137] ),
    .A2(_1163_),
    .B1(_1164_),
    .B2(\reversed_thermometer[73] ),
    .C1(_1166_),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _2949_ (.A(_1160_),
    .B(_1161_),
    .C(\reversed_thermometer[200] ),
    .X(_1167_));
 sky130_fd_sc_hd__a221o_1 _2950_ (.A1(\reversed_thermometer[136] ),
    .A2(_1163_),
    .B1(_1164_),
    .B2(\reversed_thermometer[72] ),
    .C1(_1167_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _2951_ (.A(_1160_),
    .B(_1161_),
    .C(\reversed_thermometer[199] ),
    .X(_1168_));
 sky130_fd_sc_hd__a221o_1 _2952_ (.A1(\reversed_thermometer[135] ),
    .A2(_1163_),
    .B1(_1164_),
    .B2(\reversed_thermometer[71] ),
    .C1(_1168_),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_2 _2953_ (.A(_0668_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_2 _2954_ (.A(_0671_),
    .X(_1170_));
 sky130_fd_sc_hd__and3_1 _2955_ (.A(_1169_),
    .B(_1170_),
    .C(\reversed_thermometer[198] ),
    .X(_1171_));
 sky130_fd_sc_hd__a221o_1 _2956_ (.A1(\reversed_thermometer[134] ),
    .A2(_1163_),
    .B1(_1164_),
    .B2(\reversed_thermometer[70] ),
    .C1(_1171_),
    .X(_0220_));
 sky130_fd_sc_hd__buf_2 _2957_ (.A(_0718_),
    .X(_1172_));
 sky130_fd_sc_hd__buf_2 _2958_ (.A(_0721_),
    .X(_1173_));
 sky130_fd_sc_hd__and3_1 _2959_ (.A(_1169_),
    .B(_1170_),
    .C(\reversed_thermometer[197] ),
    .X(_1174_));
 sky130_fd_sc_hd__a221o_1 _2960_ (.A1(\reversed_thermometer[133] ),
    .A2(_1172_),
    .B1(_1173_),
    .B2(\reversed_thermometer[69] ),
    .C1(_1174_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _2961_ (.A(_1169_),
    .B(_1170_),
    .C(\reversed_thermometer[196] ),
    .X(_1175_));
 sky130_fd_sc_hd__a221o_1 _2962_ (.A1(\reversed_thermometer[132] ),
    .A2(_1172_),
    .B1(_1173_),
    .B2(\reversed_thermometer[68] ),
    .C1(_1175_),
    .X(_0222_));
 sky130_fd_sc_hd__and3_1 _2963_ (.A(_1169_),
    .B(_1170_),
    .C(\reversed_thermometer[195] ),
    .X(_1176_));
 sky130_fd_sc_hd__a221o_1 _2964_ (.A1(\reversed_thermometer[131] ),
    .A2(_1172_),
    .B1(_1173_),
    .B2(\reversed_thermometer[67] ),
    .C1(_1176_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _2965_ (.A(_1169_),
    .B(_1170_),
    .C(\reversed_thermometer[194] ),
    .X(_1177_));
 sky130_fd_sc_hd__a221o_1 _2966_ (.A1(\reversed_thermometer[130] ),
    .A2(_1172_),
    .B1(_1173_),
    .B2(\reversed_thermometer[66] ),
    .C1(_1177_),
    .X(_0224_));
 sky130_fd_sc_hd__and3_1 _2967_ (.A(_0684_),
    .B(_0686_),
    .C(\reversed_thermometer[193] ),
    .X(_1178_));
 sky130_fd_sc_hd__a221o_1 _2968_ (.A1(\reversed_thermometer[129] ),
    .A2(_1172_),
    .B1(_1173_),
    .B2(\reversed_thermometer[65] ),
    .C1(_1178_),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _2969_ (.A(_0684_),
    .B(_0686_),
    .C(\reversed_thermometer[192] ),
    .X(_1179_));
 sky130_fd_sc_hd__a221o_1 _2970_ (.A1(\reversed_thermometer[128] ),
    .A2(_0675_),
    .B1(_0678_),
    .B2(\reversed_thermometer[64] ),
    .C1(_1179_),
    .X(_0226_));
 sky130_fd_sc_hd__xnor2_1 _2971_ (.A(\lfsr_q[1] ),
    .B(\lfsr_q[0] ),
    .Y(_1180_));
 sky130_fd_sc_hd__xnor2_1 _2972_ (.A(\lfsr_q[4] ),
    .B(_1180_),
    .Y(_0000_));
 sky130_fd_sc_hd__conb_1 _2973_ (.LO(_0319_));
 sky130_fd_sc_hd__buf_2 _2974_ (.A(net3),
    .X(net272));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(_0228_),
    .A1(\reversed_thermometer[255] ),
    .S(net279),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_0229_),
    .A1(\reversed_thermometer[254] ),
    .S(_0227_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_2 _2977_ (.A0(_0230_),
    .A1(\reversed_thermometer[253] ),
    .S(_0227_),
    .X(_1537_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(_0231_),
    .A1(\reversed_thermometer[252] ),
    .S(_0227_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(_0232_),
    .A1(\reversed_thermometer[251] ),
    .S(net285),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(_0233_),
    .A1(\reversed_thermometer[250] ),
    .S(net285),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_2 _2981_ (.A0(_0234_),
    .A1(\reversed_thermometer[249] ),
    .S(net286),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(_0235_),
    .A1(\reversed_thermometer[248] ),
    .S(net285),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_0236_),
    .A1(\reversed_thermometer[247] ),
    .S(net286),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(_0237_),
    .A1(\reversed_thermometer[246] ),
    .S(net285),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_2 _2985_ (.A0(_0238_),
    .A1(\reversed_thermometer[245] ),
    .S(net286),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(_0239_),
    .A1(\reversed_thermometer[244] ),
    .S(net286),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(_0240_),
    .A1(\reversed_thermometer[243] ),
    .S(net273),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(_0241_),
    .A1(\reversed_thermometer[242] ),
    .S(net273),
    .X(_1403_));
 sky130_fd_sc_hd__mux2_2 _2989_ (.A0(_0242_),
    .A1(\reversed_thermometer[241] ),
    .S(net286),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_2 _2990_ (.A0(_0243_),
    .A1(\reversed_thermometer[240] ),
    .S(net284),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_2 _2991_ (.A0(_0244_),
    .A1(\reversed_thermometer[239] ),
    .S(net284),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_2 _2992_ (.A0(_0245_),
    .A1(\reversed_thermometer[238] ),
    .S(net273),
    .X(_1447_));
 sky130_fd_sc_hd__mux2_2 _2993_ (.A0(_0246_),
    .A1(\reversed_thermometer[237] ),
    .S(net284),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(_0247_),
    .A1(\reversed_thermometer[236] ),
    .S(net284),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_2 _2995_ (.A0(_0248_),
    .A1(\reversed_thermometer[235] ),
    .S(net273),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_2 _2996_ (.A0(_0249_),
    .A1(\reversed_thermometer[234] ),
    .S(net273),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(_0250_),
    .A1(\reversed_thermometer[233] ),
    .S(net282),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(_0251_),
    .A1(\reversed_thermometer[232] ),
    .S(net284),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_2 _2999_ (.A0(_0252_),
    .A1(\reversed_thermometer[231] ),
    .S(net280),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_2 _3000_ (.A0(_0253_),
    .A1(\reversed_thermometer[230] ),
    .S(net280),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_4 _3001_ (.A0(_0254_),
    .A1(\reversed_thermometer[229] ),
    .S(net280),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(_0255_),
    .A1(\reversed_thermometer[228] ),
    .S(net280),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_2 _3003_ (.A0(_0256_),
    .A1(\reversed_thermometer[227] ),
    .S(net280),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_2 _3004_ (.A0(_0257_),
    .A1(\reversed_thermometer[226] ),
    .S(net280),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_2 _3005_ (.A0(_0258_),
    .A1(\reversed_thermometer[225] ),
    .S(net281),
    .X(_1538_));
 sky130_fd_sc_hd__mux2_2 _3006_ (.A0(_0259_),
    .A1(\reversed_thermometer[224] ),
    .S(net281),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_2 _3007_ (.A0(_0003_),
    .A1(\reversed_thermometer[223] ),
    .S(net281),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_2 _3008_ (.A0(_0004_),
    .A1(\reversed_thermometer[222] ),
    .S(net281),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(_0005_),
    .A1(\reversed_thermometer[221] ),
    .S(net281),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(_0006_),
    .A1(\reversed_thermometer[220] ),
    .S(_0227_),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(_0007_),
    .A1(\reversed_thermometer[219] ),
    .S(net279),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_2 _3012_ (.A0(_0008_),
    .A1(\reversed_thermometer[218] ),
    .S(net279),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_2 _3013_ (.A0(_0009_),
    .A1(\reversed_thermometer[217] ),
    .S(net279),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_2 _3014_ (.A0(_0010_),
    .A1(\reversed_thermometer[216] ),
    .S(net278),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(_0011_),
    .A1(\reversed_thermometer[215] ),
    .S(net278),
    .X(_1549_));
 sky130_fd_sc_hd__mux2_2 _3016_ (.A0(_0012_),
    .A1(\reversed_thermometer[214] ),
    .S(net278),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _3017_ (.A0(_0013_),
    .A1(\reversed_thermometer[213] ),
    .S(net278),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_4 _3018_ (.A0(_0014_),
    .A1(\reversed_thermometer[212] ),
    .S(net276),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_2 _3019_ (.A0(_0015_),
    .A1(\reversed_thermometer[211] ),
    .S(net276),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(_0016_),
    .A1(\reversed_thermometer[210] ),
    .S(net276),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_2 _3021_ (.A0(_0017_),
    .A1(\reversed_thermometer[209] ),
    .S(net277),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_2 _3022_ (.A0(_0018_),
    .A1(\reversed_thermometer[208] ),
    .S(net276),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(_0019_),
    .A1(\reversed_thermometer[207] ),
    .S(net277),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(_0020_),
    .A1(\reversed_thermometer[206] ),
    .S(net276),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_2 _3025_ (.A0(_0021_),
    .A1(\reversed_thermometer[205] ),
    .S(net275),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(_0022_),
    .A1(\reversed_thermometer[204] ),
    .S(net275),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(_0023_),
    .A1(\reversed_thermometer[203] ),
    .S(net275),
    .X(_1562_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(_0024_),
    .A1(\reversed_thermometer[202] ),
    .S(net275),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_4 _3029_ (.A0(_0025_),
    .A1(\reversed_thermometer[201] ),
    .S(net275),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_2 _3030_ (.A0(_0026_),
    .A1(\reversed_thermometer[200] ),
    .S(net277),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(_0027_),
    .A1(\reversed_thermometer[199] ),
    .S(net274),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_4 _3032_ (.A0(_0028_),
    .A1(\reversed_thermometer[198] ),
    .S(net274),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_2 _3033_ (.A0(_0029_),
    .A1(\reversed_thermometer[197] ),
    .S(net274),
    .X(_1568_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(_0030_),
    .A1(\reversed_thermometer[196] ),
    .S(net274),
    .X(_1569_));
 sky130_fd_sc_hd__mux2_1 _3035_ (.A0(_0031_),
    .A1(\reversed_thermometer[195] ),
    .S(net283),
    .X(_1571_));
 sky130_fd_sc_hd__mux2_2 _3036_ (.A0(_0032_),
    .A1(\reversed_thermometer[194] ),
    .S(net283),
    .X(_1572_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(_0033_),
    .A1(\reversed_thermometer[193] ),
    .S(net283),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(_0034_),
    .A1(\reversed_thermometer[192] ),
    .S(net283),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(_0035_),
    .A1(\reversed_thermometer[191] ),
    .S(net279),
    .X(_1575_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(_0036_),
    .A1(\reversed_thermometer[190] ),
    .S(_0227_),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_2 _3041_ (.A0(_0037_),
    .A1(\reversed_thermometer[189] ),
    .S(_0227_),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(_0038_),
    .A1(\reversed_thermometer[188] ),
    .S(net285),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(_0039_),
    .A1(\reversed_thermometer[187] ),
    .S(net285),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_2 _3044_ (.A0(_0040_),
    .A1(\reversed_thermometer[186] ),
    .S(net285),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_2 _3045_ (.A0(_0041_),
    .A1(\reversed_thermometer[185] ),
    .S(net285),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(_0042_),
    .A1(\reversed_thermometer[184] ),
    .S(net286),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(_0043_),
    .A1(\reversed_thermometer[183] ),
    .S(net285),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(_0044_),
    .A1(\reversed_thermometer[182] ),
    .S(net285),
    .X(_1585_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(_0045_),
    .A1(\reversed_thermometer[181] ),
    .S(net285),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_2 _3050_ (.A0(_0046_),
    .A1(\reversed_thermometer[180] ),
    .S(net283),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(_0047_),
    .A1(\reversed_thermometer[179] ),
    .S(net273),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_0048_),
    .A1(\reversed_thermometer[178] ),
    .S(net273),
    .X(_1589_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(_0049_),
    .A1(\reversed_thermometer[177] ),
    .S(net283),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_2 _3054_ (.A0(_0050_),
    .A1(\reversed_thermometer[176] ),
    .S(net286),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_2 _3055_ (.A0(_0051_),
    .A1(\reversed_thermometer[175] ),
    .S(net283),
    .X(_1593_));
 sky130_fd_sc_hd__mux2_2 _3056_ (.A0(_0052_),
    .A1(\reversed_thermometer[174] ),
    .S(net273),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(_0053_),
    .A1(\reversed_thermometer[173] ),
    .S(net273),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_2 _3058_ (.A0(_0054_),
    .A1(\reversed_thermometer[172] ),
    .S(net273),
    .X(_1596_));
 sky130_fd_sc_hd__mux2_2 _3059_ (.A0(_0055_),
    .A1(\reversed_thermometer[171] ),
    .S(net273),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_2 _3060_ (.A0(_0056_),
    .A1(\reversed_thermometer[170] ),
    .S(net282),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_0057_),
    .A1(\reversed_thermometer[169] ),
    .S(net282),
    .X(_1599_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(_0058_),
    .A1(\reversed_thermometer[168] ),
    .S(net284),
    .X(_1600_));
 sky130_fd_sc_hd__mux2_2 _3063_ (.A0(_0059_),
    .A1(\reversed_thermometer[167] ),
    .S(net282),
    .X(_1601_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(_0060_),
    .A1(\reversed_thermometer[166] ),
    .S(net280),
    .X(_1602_));
 sky130_fd_sc_hd__mux2_2 _3065_ (.A0(_0061_),
    .A1(\reversed_thermometer[165] ),
    .S(net280),
    .X(_1604_));
 sky130_fd_sc_hd__mux2_2 _3066_ (.A0(_0062_),
    .A1(\reversed_thermometer[164] ),
    .S(net280),
    .X(_1605_));
 sky130_fd_sc_hd__mux2_2 _3067_ (.A0(_0063_),
    .A1(\reversed_thermometer[163] ),
    .S(net282),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(_0064_),
    .A1(\reversed_thermometer[162] ),
    .S(net280),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_2 _3069_ (.A0(_0065_),
    .A1(\reversed_thermometer[161] ),
    .S(net282),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_2 _3070_ (.A0(_0066_),
    .A1(\reversed_thermometer[160] ),
    .S(net281),
    .X(_1609_));
 sky130_fd_sc_hd__mux2_2 _3071_ (.A0(_0067_),
    .A1(\reversed_thermometer[159] ),
    .S(net281),
    .X(_1610_));
 sky130_fd_sc_hd__mux2_2 _3072_ (.A0(_0068_),
    .A1(\reversed_thermometer[158] ),
    .S(net281),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(_0069_),
    .A1(\reversed_thermometer[157] ),
    .S(net279),
    .X(_1612_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(_0070_),
    .A1(\reversed_thermometer[156] ),
    .S(net279),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(_0071_),
    .A1(\reversed_thermometer[155] ),
    .S(net279),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_2 _3076_ (.A0(_0072_),
    .A1(\reversed_thermometer[154] ),
    .S(net279),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(_0073_),
    .A1(\reversed_thermometer[153] ),
    .S(net279),
    .X(_1362_));
 sky130_fd_sc_hd__mux2_1 _3078_ (.A0(_0074_),
    .A1(\reversed_thermometer[152] ),
    .S(net278),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(_0075_),
    .A1(\reversed_thermometer[151] ),
    .S(net278),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_4 _3080_ (.A0(_0076_),
    .A1(\reversed_thermometer[150] ),
    .S(net278),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_2 _3081_ (.A0(_0077_),
    .A1(\reversed_thermometer[149] ),
    .S(net278),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_2 _3082_ (.A0(_0078_),
    .A1(\reversed_thermometer[148] ),
    .S(net276),
    .X(_1367_));
 sky130_fd_sc_hd__mux2_2 _3083_ (.A0(_0079_),
    .A1(\reversed_thermometer[147] ),
    .S(net276),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_2 _3084_ (.A0(_0080_),
    .A1(\reversed_thermometer[146] ),
    .S(net277),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_2 _3085_ (.A0(_0081_),
    .A1(\reversed_thermometer[145] ),
    .S(net277),
    .X(_1371_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(_0082_),
    .A1(\reversed_thermometer[144] ),
    .S(net276),
    .X(_1372_));
 sky130_fd_sc_hd__mux2_4 _3087_ (.A0(_0083_),
    .A1(\reversed_thermometer[143] ),
    .S(net277),
    .X(_1373_));
 sky130_fd_sc_hd__mux2_2 _3088_ (.A0(_0084_),
    .A1(\reversed_thermometer[142] ),
    .S(net276),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(_0085_),
    .A1(\reversed_thermometer[141] ),
    .S(net277),
    .X(_1375_));
 sky130_fd_sc_hd__mux2_4 _3090_ (.A0(_0086_),
    .A1(\reversed_thermometer[140] ),
    .S(net275),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(_0087_),
    .A1(\reversed_thermometer[139] ),
    .S(net275),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_4 _3092_ (.A0(_0088_),
    .A1(\reversed_thermometer[138] ),
    .S(net275),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(_0089_),
    .A1(\reversed_thermometer[137] ),
    .S(net275),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(_0090_),
    .A1(\reversed_thermometer[136] ),
    .S(net277),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_2 _3095_ (.A0(_0091_),
    .A1(\reversed_thermometer[135] ),
    .S(net274),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(_0092_),
    .A1(\reversed_thermometer[134] ),
    .S(net274),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(_0093_),
    .A1(\reversed_thermometer[133] ),
    .S(net274),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_4 _3098_ (.A0(_0094_),
    .A1(\reversed_thermometer[132] ),
    .S(net274),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_2 _3099_ (.A0(_0095_),
    .A1(\reversed_thermometer[131] ),
    .S(net283),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_2 _3100_ (.A0(_0096_),
    .A1(\reversed_thermometer[130] ),
    .S(net283),
    .X(_1387_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_0097_),
    .A1(\reversed_thermometer[129] ),
    .S(net283),
    .X(_1388_));
 sky130_fd_sc_hd__mux2_1 _3102_ (.A0(_0098_),
    .A1(\reversed_thermometer[128] ),
    .S(net283),
    .X(_1389_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_0099_),
    .A1(\reversed_thermometer[127] ),
    .S(net279),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(_0100_),
    .A1(\reversed_thermometer[126] ),
    .S(_0227_),
    .X(_1391_));
 sky130_fd_sc_hd__mux2_2 _3105_ (.A0(_0101_),
    .A1(\reversed_thermometer[125] ),
    .S(net285),
    .X(_1393_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(_0102_),
    .A1(\reversed_thermometer[124] ),
    .S(_0227_),
    .X(_1394_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_0103_),
    .A1(\reversed_thermometer[123] ),
    .S(net285),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_2 _3108_ (.A0(_0104_),
    .A1(\reversed_thermometer[122] ),
    .S(net286),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(_0105_),
    .A1(\reversed_thermometer[121] ),
    .S(net285),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_2 _3110_ (.A0(_0106_),
    .A1(\reversed_thermometer[120] ),
    .S(net286),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(_0107_),
    .A1(\reversed_thermometer[119] ),
    .S(net286),
    .X(_1399_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(_0108_),
    .A1(\reversed_thermometer[118] ),
    .S(net286),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_2 _3113_ (.A0(_0109_),
    .A1(\reversed_thermometer[117] ),
    .S(net286),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(_0110_),
    .A1(\reversed_thermometer[116] ),
    .S(net286),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(_0111_),
    .A1(\reversed_thermometer[115] ),
    .S(net273),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_2 _3116_ (.A0(_0112_),
    .A1(\reversed_thermometer[114] ),
    .S(net273),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_2 _3117_ (.A0(_0113_),
    .A1(\reversed_thermometer[113] ),
    .S(net286),
    .X(_1406_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(_0114_),
    .A1(\reversed_thermometer[112] ),
    .S(net284),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(_0115_),
    .A1(\reversed_thermometer[111] ),
    .S(net284),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(_0116_),
    .A1(\reversed_thermometer[110] ),
    .S(net284),
    .X(_1409_));
 sky130_fd_sc_hd__mux2_2 _3121_ (.A0(_0117_),
    .A1(\reversed_thermometer[109] ),
    .S(net284),
    .X(_1410_));
 sky130_fd_sc_hd__mux2_2 _3122_ (.A0(_0118_),
    .A1(\reversed_thermometer[108] ),
    .S(net284),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(_0119_),
    .A1(\reversed_thermometer[107] ),
    .S(net284),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_2 _3124_ (.A0(_0120_),
    .A1(\reversed_thermometer[106] ),
    .S(net284),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(_0121_),
    .A1(\reversed_thermometer[105] ),
    .S(net282),
    .X(_1415_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(_0122_),
    .A1(\reversed_thermometer[104] ),
    .S(net284),
    .X(_1416_));
 sky130_fd_sc_hd__mux2_2 _3127_ (.A0(_0123_),
    .A1(\reversed_thermometer[103] ),
    .S(net282),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_2 _3128_ (.A0(_0124_),
    .A1(\reversed_thermometer[102] ),
    .S(net280),
    .X(_1418_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(_0125_),
    .A1(\reversed_thermometer[101] ),
    .S(net280),
    .X(_1419_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(_0126_),
    .A1(\reversed_thermometer[100] ),
    .S(net280),
    .X(_1420_));
 sky130_fd_sc_hd__mux2_2 _3131_ (.A0(_0127_),
    .A1(\reversed_thermometer[99] ),
    .S(net282),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(_0128_),
    .A1(\reversed_thermometer[98] ),
    .S(net280),
    .X(_1422_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(_0129_),
    .A1(\reversed_thermometer[97] ),
    .S(net282),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(_0130_),
    .A1(\reversed_thermometer[96] ),
    .S(net281),
    .X(_1424_));
 sky130_fd_sc_hd__mux2_2 _3135_ (.A0(_0131_),
    .A1(\reversed_thermometer[95] ),
    .S(net281),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_2 _3136_ (.A0(_0132_),
    .A1(\reversed_thermometer[94] ),
    .S(net281),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_2 _3137_ (.A0(_0133_),
    .A1(\reversed_thermometer[93] ),
    .S(net279),
    .X(_1428_));
 sky130_fd_sc_hd__mux2_2 _3138_ (.A0(_0134_),
    .A1(\reversed_thermometer[92] ),
    .S(_0227_),
    .X(_1429_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(_0135_),
    .A1(\reversed_thermometer[91] ),
    .S(_0227_),
    .X(_1430_));
 sky130_fd_sc_hd__mux2_2 _3140_ (.A0(_0136_),
    .A1(\reversed_thermometer[90] ),
    .S(net278),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_2 _3141_ (.A0(_0137_),
    .A1(\reversed_thermometer[89] ),
    .S(net279),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_2 _3142_ (.A0(_0138_),
    .A1(\reversed_thermometer[88] ),
    .S(net278),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_2 _3143_ (.A0(_0139_),
    .A1(\reversed_thermometer[87] ),
    .S(net278),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_2 _3144_ (.A0(_0140_),
    .A1(\reversed_thermometer[86] ),
    .S(net278),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(_0141_),
    .A1(\reversed_thermometer[85] ),
    .S(net278),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(_0142_),
    .A1(\reversed_thermometer[84] ),
    .S(net276),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(_0143_),
    .A1(\reversed_thermometer[83] ),
    .S(net276),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_2 _3148_ (.A0(_0144_),
    .A1(\reversed_thermometer[82] ),
    .S(net277),
    .X(_1440_));
 sky130_fd_sc_hd__mux2_2 _3149_ (.A0(_0145_),
    .A1(\reversed_thermometer[81] ),
    .S(net277),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(_0146_),
    .A1(\reversed_thermometer[80] ),
    .S(net276),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_1 _3151_ (.A0(_0147_),
    .A1(\reversed_thermometer[79] ),
    .S(net277),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(_0148_),
    .A1(\reversed_thermometer[78] ),
    .S(net276),
    .X(_1444_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(_0149_),
    .A1(\reversed_thermometer[77] ),
    .S(net276),
    .X(_1445_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(_0150_),
    .A1(\reversed_thermometer[76] ),
    .S(net275),
    .X(_1446_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(_0151_),
    .A1(\reversed_thermometer[75] ),
    .S(net275),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(_0152_),
    .A1(\reversed_thermometer[74] ),
    .S(net275),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(_0153_),
    .A1(\reversed_thermometer[73] ),
    .S(net275),
    .X(_1450_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(_0154_),
    .A1(\reversed_thermometer[72] ),
    .S(net277),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_2 _3159_ (.A0(_0155_),
    .A1(\reversed_thermometer[71] ),
    .S(net274),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(_0156_),
    .A1(\reversed_thermometer[70] ),
    .S(net274),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _3161_ (.A0(_0157_),
    .A1(\reversed_thermometer[69] ),
    .S(net274),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(_0158_),
    .A1(\reversed_thermometer[68] ),
    .S(net274),
    .X(_1455_));
 sky130_fd_sc_hd__mux2_2 _3163_ (.A0(_0159_),
    .A1(\reversed_thermometer[67] ),
    .S(net280),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(_0160_),
    .A1(\reversed_thermometer[66] ),
    .S(net280),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_2 _3165_ (.A0(_0161_),
    .A1(\reversed_thermometer[65] ),
    .S(net283),
    .X(_1459_));
 sky130_fd_sc_hd__mux2_2 _3166_ (.A0(_0162_),
    .A1(\reversed_thermometer[64] ),
    .S(net283),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(_0163_),
    .A1(\reversed_thermometer[63] ),
    .S(net279),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(_0164_),
    .A1(\reversed_thermometer[62] ),
    .S(_0227_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_0165_),
    .A1(\reversed_thermometer[61] ),
    .S(net285),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_2 _3170_ (.A0(_0166_),
    .A1(\reversed_thermometer[60] ),
    .S(net285),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(_0167_),
    .A1(\reversed_thermometer[59] ),
    .S(net285),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_2 _3172_ (.A0(_0168_),
    .A1(\reversed_thermometer[58] ),
    .S(net285),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(_0169_),
    .A1(\reversed_thermometer[57] ),
    .S(net285),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _3174_ (.A0(_0170_),
    .A1(\reversed_thermometer[56] ),
    .S(net286),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(_0171_),
    .A1(\reversed_thermometer[55] ),
    .S(net285),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _3176_ (.A0(_0172_),
    .A1(\reversed_thermometer[54] ),
    .S(net286),
    .X(_1472_));
 sky130_fd_sc_hd__mux2_2 _3177_ (.A0(_0173_),
    .A1(\reversed_thermometer[53] ),
    .S(net286),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_2 _3178_ (.A0(_0174_),
    .A1(\reversed_thermometer[52] ),
    .S(net283),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(_0175_),
    .A1(\reversed_thermometer[51] ),
    .S(net273),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_2 _3180_ (.A0(_0176_),
    .A1(\reversed_thermometer[50] ),
    .S(net273),
    .X(_1476_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(_0177_),
    .A1(\reversed_thermometer[49] ),
    .S(net286),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(_0178_),
    .A1(\reversed_thermometer[48] ),
    .S(net284),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(_0179_),
    .A1(\reversed_thermometer[47] ),
    .S(net273),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(_0180_),
    .A1(\reversed_thermometer[46] ),
    .S(net273),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(_0181_),
    .A1(\reversed_thermometer[45] ),
    .S(net273),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(_0182_),
    .A1(\reversed_thermometer[44] ),
    .S(net273),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_2 _3187_ (.A0(_0183_),
    .A1(\reversed_thermometer[43] ),
    .S(net273),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_2 _3188_ (.A0(_0184_),
    .A1(\reversed_thermometer[42] ),
    .S(net273),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(_0185_),
    .A1(\reversed_thermometer[41] ),
    .S(net282),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_2 _3190_ (.A0(_0186_),
    .A1(\reversed_thermometer[40] ),
    .S(net284),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(_0187_),
    .A1(\reversed_thermometer[39] ),
    .S(net282),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(_0188_),
    .A1(\reversed_thermometer[38] ),
    .S(net280),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_2 _3193_ (.A0(_0189_),
    .A1(\reversed_thermometer[37] ),
    .S(net280),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(_0190_),
    .A1(\reversed_thermometer[36] ),
    .S(net280),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(_0191_),
    .A1(\reversed_thermometer[35] ),
    .S(net282),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_2 _3196_ (.A0(_0192_),
    .A1(\reversed_thermometer[34] ),
    .S(net280),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_2 _3197_ (.A0(_0193_),
    .A1(\reversed_thermometer[33] ),
    .S(net281),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(_0194_),
    .A1(\reversed_thermometer[32] ),
    .S(net281),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_2 _3199_ (.A0(_0195_),
    .A1(\reversed_thermometer[31] ),
    .S(net281),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(_0196_),
    .A1(\reversed_thermometer[30] ),
    .S(net279),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_2 _3201_ (.A0(_0197_),
    .A1(\reversed_thermometer[29] ),
    .S(net279),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(_0198_),
    .A1(\reversed_thermometer[28] ),
    .S(_0227_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_2 _3203_ (.A0(_0199_),
    .A1(\reversed_thermometer[27] ),
    .S(net279),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_2 _3204_ (.A0(_0200_),
    .A1(\reversed_thermometer[26] ),
    .S(net279),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_4 _3205_ (.A0(_0201_),
    .A1(\reversed_thermometer[25] ),
    .S(net279),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_2 _3206_ (.A0(_0202_),
    .A1(\reversed_thermometer[24] ),
    .S(net278),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_2 _3207_ (.A0(_0203_),
    .A1(\reversed_thermometer[23] ),
    .S(net278),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(_0204_),
    .A1(\reversed_thermometer[22] ),
    .S(net278),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(_0205_),
    .A1(\reversed_thermometer[21] ),
    .S(net278),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_4 _3210_ (.A0(_0206_),
    .A1(\reversed_thermometer[20] ),
    .S(net276),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_4 _3211_ (.A0(_0207_),
    .A1(\reversed_thermometer[19] ),
    .S(net276),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_2 _3212_ (.A0(_0208_),
    .A1(\reversed_thermometer[18] ),
    .S(net277),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_2 _3213_ (.A0(_0209_),
    .A1(\reversed_thermometer[17] ),
    .S(net277),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(_0210_),
    .A1(\reversed_thermometer[16] ),
    .S(net276),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_2 _3215_ (.A0(_0211_),
    .A1(\reversed_thermometer[15] ),
    .S(net277),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_4 _3216_ (.A0(_0212_),
    .A1(\reversed_thermometer[14] ),
    .S(net276),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(_0213_),
    .A1(\reversed_thermometer[13] ),
    .S(net277),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(_0214_),
    .A1(\reversed_thermometer[12] ),
    .S(net275),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_4 _3219_ (.A0(_0215_),
    .A1(\reversed_thermometer[11] ),
    .S(net275),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_4 _3220_ (.A0(_0216_),
    .A1(\reversed_thermometer[10] ),
    .S(net275),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(_0217_),
    .A1(\reversed_thermometer[9] ),
    .S(net275),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(_0218_),
    .A1(\reversed_thermometer[8] ),
    .S(net277),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(_0219_),
    .A1(\reversed_thermometer[7] ),
    .S(net274),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(_0220_),
    .A1(\reversed_thermometer[6] ),
    .S(net274),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_4 _3225_ (.A0(_0221_),
    .A1(\reversed_thermometer[5] ),
    .S(net274),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_4 _3226_ (.A0(_0222_),
    .A1(\reversed_thermometer[4] ),
    .S(net274),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_2 _3227_ (.A0(_0223_),
    .A1(\reversed_thermometer[3] ),
    .S(net280),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_2 _3228_ (.A0(_0224_),
    .A1(\reversed_thermometer[2] ),
    .S(net281),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(_0225_),
    .A1(\reversed_thermometer[1] ),
    .S(net281),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(_0226_),
    .A1(\reversed_thermometer[0] ),
    .S(net283),
    .X(_1531_));
 sky130_fd_sc_hd__dfxtp_1 _3231_ (.D(_0260_),
    .Q(\reversed_thermometer[196] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3232_ (.D(_0261_),
    .Q(\reversed_thermometer[197] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3233_ (.D(_0262_),
    .Q(\reversed_thermometer[198] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3234_ (.D(_0263_),
    .Q(\reversed_thermometer[199] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3235_ (.D(_0264_),
    .Q(\reversed_thermometer[200] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3236_ (.D(_0265_),
    .Q(\reversed_thermometer[201] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3237_ (.D(_0266_),
    .Q(\reversed_thermometer[202] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3238_ (.D(_0267_),
    .Q(\reversed_thermometer[203] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3239_ (.D(_0268_),
    .Q(\reversed_thermometer[204] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3240_ (.D(_0269_),
    .Q(\reversed_thermometer[205] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3241_ (.D(_0270_),
    .Q(\reversed_thermometer[206] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3242_ (.D(_0271_),
    .Q(\reversed_thermometer[207] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3243_ (.D(_0272_),
    .Q(\reversed_thermometer[208] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3244_ (.D(_0273_),
    .Q(\reversed_thermometer[209] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3245_ (.D(_0274_),
    .Q(\reversed_thermometer[210] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3246_ (.D(_0275_),
    .Q(\reversed_thermometer[211] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3247_ (.D(_0276_),
    .Q(\reversed_thermometer[212] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3248_ (.D(_0277_),
    .Q(\reversed_thermometer[213] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3249_ (.D(_0278_),
    .Q(\reversed_thermometer[214] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3250_ (.D(_0279_),
    .Q(\reversed_thermometer[215] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3251_ (.D(_0280_),
    .Q(\reversed_thermometer[216] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3252_ (.D(_0281_),
    .Q(\reversed_thermometer[217] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3253_ (.D(_0282_),
    .Q(\reversed_thermometer[218] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3254_ (.D(_0283_),
    .Q(\reversed_thermometer[219] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3255_ (.D(_0284_),
    .Q(\reversed_thermometer[220] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3256_ (.D(_0285_),
    .Q(\reversed_thermometer[221] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3257_ (.D(_0286_),
    .Q(\reversed_thermometer[222] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3258_ (.D(_0287_),
    .Q(\reversed_thermometer[223] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3259_ (.D(_0288_),
    .Q(\reversed_thermometer[224] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3260_ (.D(_0289_),
    .Q(\reversed_thermometer[225] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3261_ (.D(_0290_),
    .Q(\reversed_thermometer[226] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3262_ (.D(_0291_),
    .Q(\reversed_thermometer[227] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3263_ (.D(_0292_),
    .Q(\reversed_thermometer[228] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3264_ (.D(_0293_),
    .Q(\reversed_thermometer[229] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3265_ (.D(_0294_),
    .Q(\reversed_thermometer[230] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3266_ (.D(_0295_),
    .Q(\reversed_thermometer[231] ),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3267_ (.D(_0296_),
    .Q(\reversed_thermometer[232] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3268_ (.D(_0297_),
    .Q(\reversed_thermometer[233] ),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3269_ (.D(_0298_),
    .Q(\reversed_thermometer[234] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3270_ (.D(_0299_),
    .Q(\reversed_thermometer[235] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3271_ (.D(_0300_),
    .Q(\reversed_thermometer[236] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3272_ (.D(_0301_),
    .Q(\reversed_thermometer[237] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3273_ (.D(_0302_),
    .Q(\reversed_thermometer[238] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3274_ (.D(_0303_),
    .Q(\reversed_thermometer[239] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3275_ (.D(_0304_),
    .Q(\reversed_thermometer[240] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3276_ (.D(_0305_),
    .Q(\reversed_thermometer[241] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3277_ (.D(_0306_),
    .Q(\reversed_thermometer[242] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3278_ (.D(_0307_),
    .Q(\reversed_thermometer[243] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3279_ (.D(_0308_),
    .Q(\reversed_thermometer[244] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3280_ (.D(_0309_),
    .Q(\reversed_thermometer[245] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3281_ (.D(_0310_),
    .Q(\reversed_thermometer[246] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3282_ (.D(_0311_),
    .Q(\reversed_thermometer[247] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3283_ (.D(_0312_),
    .Q(\reversed_thermometer[248] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3284_ (.D(_0313_),
    .Q(\reversed_thermometer[249] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3285_ (.D(_0314_),
    .Q(\reversed_thermometer[250] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3286_ (.D(_0315_),
    .Q(\reversed_thermometer[251] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3287_ (.D(_0316_),
    .Q(\reversed_thermometer[252] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3288_ (.D(_0317_),
    .Q(\reversed_thermometer[253] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3289_ (.D(_0318_),
    .Q(\reversed_thermometer[254] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3290_ (.D(_0319_),
    .Q(\reversed_thermometer[0] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3291_ (.D(_0320_),
    .Q(\reversed_thermometer[1] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3292_ (.D(_0321_),
    .Q(\reversed_thermometer[2] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3293_ (.D(_0322_),
    .Q(\reversed_thermometer[3] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3294_ (.D(_0323_),
    .Q(\reversed_thermometer[4] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3295_ (.D(_0324_),
    .Q(\reversed_thermometer[5] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3296_ (.D(_0325_),
    .Q(\reversed_thermometer[6] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3297_ (.D(_0326_),
    .Q(\reversed_thermometer[7] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3298_ (.D(_0327_),
    .Q(\reversed_thermometer[8] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3299_ (.D(_0328_),
    .Q(\reversed_thermometer[9] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3300_ (.D(_0329_),
    .Q(\reversed_thermometer[10] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3301_ (.D(_0330_),
    .Q(\reversed_thermometer[11] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3302_ (.D(_0331_),
    .Q(\reversed_thermometer[12] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3303_ (.D(_0332_),
    .Q(\reversed_thermometer[13] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3304_ (.D(_0333_),
    .Q(\reversed_thermometer[14] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.D(_0334_),
    .Q(\reversed_thermometer[15] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.D(_0335_),
    .Q(\reversed_thermometer[16] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3307_ (.D(_0336_),
    .Q(\reversed_thermometer[17] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3308_ (.D(_0337_),
    .Q(\reversed_thermometer[18] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3309_ (.D(_0338_),
    .Q(\reversed_thermometer[19] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3310_ (.D(_0339_),
    .Q(\reversed_thermometer[20] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3311_ (.D(_0340_),
    .Q(\reversed_thermometer[21] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3312_ (.D(_0341_),
    .Q(\reversed_thermometer[22] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3313_ (.D(_0342_),
    .Q(\reversed_thermometer[23] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3314_ (.D(_0343_),
    .Q(\reversed_thermometer[24] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3315_ (.D(_0344_),
    .Q(\reversed_thermometer[25] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3316_ (.D(_0345_),
    .Q(\reversed_thermometer[26] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3317_ (.D(_0346_),
    .Q(\reversed_thermometer[27] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3318_ (.D(_0347_),
    .Q(\reversed_thermometer[28] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3319_ (.D(_0348_),
    .Q(\reversed_thermometer[29] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3320_ (.D(_0349_),
    .Q(\reversed_thermometer[30] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3321_ (.D(_0350_),
    .Q(\reversed_thermometer[31] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3322_ (.D(_0351_),
    .Q(\reversed_thermometer[32] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3323_ (.D(_0352_),
    .Q(\reversed_thermometer[33] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3324_ (.D(_0353_),
    .Q(\reversed_thermometer[34] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.D(_0354_),
    .Q(\reversed_thermometer[35] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3326_ (.D(_0355_),
    .Q(\reversed_thermometer[36] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.D(_0356_),
    .Q(\reversed_thermometer[37] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.D(_0357_),
    .Q(\reversed_thermometer[38] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.D(_0358_),
    .Q(\reversed_thermometer[39] ),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.D(_0359_),
    .Q(\reversed_thermometer[40] ),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.D(_0360_),
    .Q(\reversed_thermometer[41] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.D(_0361_),
    .Q(\reversed_thermometer[42] ),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.D(_0362_),
    .Q(\reversed_thermometer[43] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.D(_0363_),
    .Q(\reversed_thermometer[44] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.D(_0364_),
    .Q(\reversed_thermometer[45] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.D(_0365_),
    .Q(\reversed_thermometer[46] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.D(_0366_),
    .Q(\reversed_thermometer[47] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.D(_0367_),
    .Q(\reversed_thermometer[48] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.D(_0368_),
    .Q(\reversed_thermometer[49] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3340_ (.D(_0369_),
    .Q(\reversed_thermometer[50] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3341_ (.D(_0370_),
    .Q(\reversed_thermometer[51] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.D(_0371_),
    .Q(\reversed_thermometer[52] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.D(_0372_),
    .Q(\reversed_thermometer[53] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3344_ (.D(_0373_),
    .Q(\reversed_thermometer[54] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3345_ (.D(_0374_),
    .Q(\reversed_thermometer[55] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3346_ (.D(_0375_),
    .Q(\reversed_thermometer[56] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3347_ (.D(_0376_),
    .Q(\reversed_thermometer[57] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3348_ (.D(_0377_),
    .Q(\reversed_thermometer[58] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3349_ (.D(_0378_),
    .Q(\reversed_thermometer[59] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3350_ (.D(_0379_),
    .Q(\reversed_thermometer[60] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3351_ (.D(_0380_),
    .Q(\reversed_thermometer[61] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3352_ (.D(_0381_),
    .Q(\reversed_thermometer[62] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3353_ (.D(_0382_),
    .Q(\reversed_thermometer[63] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3354_ (.D(_0383_),
    .Q(\reversed_thermometer[64] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3355_ (.D(_0384_),
    .Q(\reversed_thermometer[65] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3356_ (.D(_0385_),
    .Q(\reversed_thermometer[66] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3357_ (.D(_0386_),
    .Q(\reversed_thermometer[67] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3358_ (.D(_0387_),
    .Q(\reversed_thermometer[68] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3359_ (.D(_0388_),
    .Q(\reversed_thermometer[69] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.D(_0389_),
    .Q(\reversed_thermometer[70] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.D(_0390_),
    .Q(\reversed_thermometer[71] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.D(_0391_),
    .Q(\reversed_thermometer[72] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.D(_0392_),
    .Q(\reversed_thermometer[73] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.D(_0393_),
    .Q(\reversed_thermometer[74] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.D(_0394_),
    .Q(\reversed_thermometer[75] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.D(_0395_),
    .Q(\reversed_thermometer[76] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.D(_0396_),
    .Q(\reversed_thermometer[77] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.D(_0397_),
    .Q(\reversed_thermometer[78] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.D(_0398_),
    .Q(\reversed_thermometer[79] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.D(_0399_),
    .Q(\reversed_thermometer[80] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3371_ (.D(_0400_),
    .Q(\reversed_thermometer[81] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3372_ (.D(_0401_),
    .Q(\reversed_thermometer[82] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3373_ (.D(_0402_),
    .Q(\reversed_thermometer[83] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3374_ (.D(_0403_),
    .Q(\reversed_thermometer[84] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3375_ (.D(_0404_),
    .Q(\reversed_thermometer[85] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.D(_0405_),
    .Q(\reversed_thermometer[86] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.D(_0406_),
    .Q(\reversed_thermometer[87] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.D(_0407_),
    .Q(\reversed_thermometer[88] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.D(_0408_),
    .Q(\reversed_thermometer[89] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3380_ (.D(_0409_),
    .Q(\reversed_thermometer[90] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3381_ (.D(_0410_),
    .Q(\reversed_thermometer[91] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.D(_0411_),
    .Q(\reversed_thermometer[92] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3383_ (.D(_0412_),
    .Q(\reversed_thermometer[93] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3384_ (.D(_0413_),
    .Q(\reversed_thermometer[94] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3385_ (.D(_0414_),
    .Q(\reversed_thermometer[95] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3386_ (.D(_0415_),
    .Q(\reversed_thermometer[96] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3387_ (.D(_0416_),
    .Q(\reversed_thermometer[97] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3388_ (.D(_0417_),
    .Q(\reversed_thermometer[98] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3389_ (.D(_0418_),
    .Q(\reversed_thermometer[99] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3390_ (.D(_0419_),
    .Q(\reversed_thermometer[100] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3391_ (.D(_0420_),
    .Q(\reversed_thermometer[101] ),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3392_ (.D(_0421_),
    .Q(\reversed_thermometer[102] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3393_ (.D(_0422_),
    .Q(\reversed_thermometer[103] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3394_ (.D(_0423_),
    .Q(\reversed_thermometer[104] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3395_ (.D(_0424_),
    .Q(\reversed_thermometer[105] ),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3396_ (.D(_0425_),
    .Q(\reversed_thermometer[106] ),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3397_ (.D(_0426_),
    .Q(\reversed_thermometer[107] ),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3398_ (.D(_0427_),
    .Q(\reversed_thermometer[108] ),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3399_ (.D(_0428_),
    .Q(\reversed_thermometer[109] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3400_ (.D(_0429_),
    .Q(\reversed_thermometer[110] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3401_ (.D(_0430_),
    .Q(\reversed_thermometer[111] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3402_ (.D(_0431_),
    .Q(\reversed_thermometer[112] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3403_ (.D(_0432_),
    .Q(\reversed_thermometer[113] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3404_ (.D(_0433_),
    .Q(\reversed_thermometer[114] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3405_ (.D(_0434_),
    .Q(\reversed_thermometer[115] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3406_ (.D(_0435_),
    .Q(\reversed_thermometer[116] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3407_ (.D(_0436_),
    .Q(\reversed_thermometer[117] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3408_ (.D(_0437_),
    .Q(\reversed_thermometer[118] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3409_ (.D(_0438_),
    .Q(\reversed_thermometer[119] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3410_ (.D(_0439_),
    .Q(\reversed_thermometer[120] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3411_ (.D(_0440_),
    .Q(\reversed_thermometer[121] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3412_ (.D(_0441_),
    .Q(\reversed_thermometer[122] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3413_ (.D(_0442_),
    .Q(\reversed_thermometer[123] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3414_ (.D(_0443_),
    .Q(\reversed_thermometer[124] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3415_ (.D(_0444_),
    .Q(\reversed_thermometer[125] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3416_ (.D(_0445_),
    .Q(\reversed_thermometer[126] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3417_ (.D(_0446_),
    .Q(\reversed_thermometer[127] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3418_ (.D(_0447_),
    .Q(\reversed_thermometer[128] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3419_ (.D(_0448_),
    .Q(\reversed_thermometer[129] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3420_ (.D(_0449_),
    .Q(\reversed_thermometer[130] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3421_ (.D(_0450_),
    .Q(\reversed_thermometer[131] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3422_ (.D(_0451_),
    .Q(\reversed_thermometer[132] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3423_ (.D(_0452_),
    .Q(\reversed_thermometer[133] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3424_ (.D(_0453_),
    .Q(\reversed_thermometer[134] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3425_ (.D(_0454_),
    .Q(\reversed_thermometer[135] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3426_ (.D(_0455_),
    .Q(\reversed_thermometer[136] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3427_ (.D(_0456_),
    .Q(\reversed_thermometer[137] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3428_ (.D(_0457_),
    .Q(\reversed_thermometer[138] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3429_ (.D(_0458_),
    .Q(\reversed_thermometer[139] ),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3430_ (.D(_0459_),
    .Q(\reversed_thermometer[140] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3431_ (.D(_0460_),
    .Q(\reversed_thermometer[141] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3432_ (.D(_0461_),
    .Q(\reversed_thermometer[142] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3433_ (.D(_0462_),
    .Q(\reversed_thermometer[143] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3434_ (.D(_0463_),
    .Q(\reversed_thermometer[144] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3435_ (.D(_0464_),
    .Q(\reversed_thermometer[145] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3436_ (.D(_0465_),
    .Q(\reversed_thermometer[146] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3437_ (.D(_0466_),
    .Q(\reversed_thermometer[147] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3438_ (.D(_0467_),
    .Q(\reversed_thermometer[148] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3439_ (.D(_0468_),
    .Q(\reversed_thermometer[149] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3440_ (.D(_0469_),
    .Q(\reversed_thermometer[150] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3441_ (.D(_0470_),
    .Q(\reversed_thermometer[151] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3442_ (.D(_0471_),
    .Q(\reversed_thermometer[152] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3443_ (.D(_0472_),
    .Q(\reversed_thermometer[153] ),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3444_ (.D(_0473_),
    .Q(\reversed_thermometer[154] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3445_ (.D(_0474_),
    .Q(\reversed_thermometer[155] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3446_ (.D(_0475_),
    .Q(\reversed_thermometer[156] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3447_ (.D(_0476_),
    .Q(\reversed_thermometer[157] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3448_ (.D(_0477_),
    .Q(\reversed_thermometer[158] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3449_ (.D(_0478_),
    .Q(\reversed_thermometer[159] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3450_ (.D(_0479_),
    .Q(\reversed_thermometer[160] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3451_ (.D(_0480_),
    .Q(\reversed_thermometer[161] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3452_ (.D(_0481_),
    .Q(\reversed_thermometer[162] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3453_ (.D(_0482_),
    .Q(\reversed_thermometer[163] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3454_ (.D(_0483_),
    .Q(\reversed_thermometer[164] ),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3455_ (.D(_0484_),
    .Q(\reversed_thermometer[165] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3456_ (.D(_0485_),
    .Q(\reversed_thermometer[166] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3457_ (.D(_0486_),
    .Q(\reversed_thermometer[167] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3458_ (.D(_0487_),
    .Q(\reversed_thermometer[168] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.D(_0488_),
    .Q(\reversed_thermometer[169] ),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.D(_0489_),
    .Q(\reversed_thermometer[170] ),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.D(_0490_),
    .Q(\reversed_thermometer[171] ),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.D(_0491_),
    .Q(\reversed_thermometer[172] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.D(_0492_),
    .Q(\reversed_thermometer[173] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.D(_0493_),
    .Q(\reversed_thermometer[174] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.D(_0494_),
    .Q(\reversed_thermometer[175] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.D(_0495_),
    .Q(\reversed_thermometer[176] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3467_ (.D(_0496_),
    .Q(\reversed_thermometer[177] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.D(_0497_),
    .Q(\reversed_thermometer[178] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3469_ (.D(_0498_),
    .Q(\reversed_thermometer[179] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3470_ (.D(_0499_),
    .Q(\reversed_thermometer[180] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3471_ (.D(_0500_),
    .Q(\reversed_thermometer[181] ),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.D(_0501_),
    .Q(\reversed_thermometer[182] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.D(_0502_),
    .Q(\reversed_thermometer[183] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.D(_0503_),
    .Q(\reversed_thermometer[184] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.D(_0504_),
    .Q(\reversed_thermometer[185] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.D(_0505_),
    .Q(\reversed_thermometer[186] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.D(_0506_),
    .Q(\reversed_thermometer[187] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.D(_0507_),
    .Q(\reversed_thermometer[188] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.D(_0508_),
    .Q(\reversed_thermometer[189] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.D(_0509_),
    .Q(\reversed_thermometer[190] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.D(_0510_),
    .Q(\reversed_thermometer[191] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.D(_0511_),
    .Q(\reversed_thermometer[192] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.D(_0512_),
    .Q(\reversed_thermometer[193] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.D(_0513_),
    .Q(\reversed_thermometer[194] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.D(_0514_),
    .Q(\reversed_thermometer[195] ),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.D(_1359_),
    .Q(net269),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.D(_1470_),
    .Q(net223),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.D(_1537_),
    .Q(net132),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.D(_1548_),
    .Q(net133),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.D(_1559_),
    .Q(net27),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.D(_1570_),
    .Q(net71),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.D(_1581_),
    .Q(net267),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.D(_1592_),
    .Q(net94),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.D(_1603_),
    .Q(net136),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.D(_1614_),
    .Q(net58),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.D(_1370_),
    .Q(net211),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.D(_1381_),
    .Q(net74),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.D(_1392_),
    .Q(net65),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.D(_1403_),
    .Q(net162),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.D(_1414_),
    .Q(net53),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.D(_1425_),
    .Q(net23),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.D(_1436_),
    .Q(net141),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.D(_1447_),
    .Q(net21),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.D(_1458_),
    .Q(net119),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.D(_1469_),
    .Q(net150),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.D(_1481_),
    .Q(net91),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.D(_1492_),
    .Q(net95),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.D(_1503_),
    .Q(net234),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.D(_1514_),
    .Q(net110),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.D(_1525_),
    .Q(net271),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.D(_1532_),
    .Q(net157),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.D(_1533_),
    .Q(net121),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.D(_1534_),
    .Q(net124),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.D(_1535_),
    .Q(net241),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.D(_1536_),
    .Q(net68),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.D(_1538_),
    .Q(net82),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.D(_1539_),
    .Q(net89),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.D(_1540_),
    .Q(net92),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.D(_1541_),
    .Q(net72),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.D(_1542_),
    .Q(net205),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.D(_1543_),
    .Q(net153),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.D(_1544_),
    .Q(net225),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.D(_1545_),
    .Q(net98),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.D(_1546_),
    .Q(net252),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.D(_1547_),
    .Q(net172),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.D(_1549_),
    .Q(net215),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.D(_1550_),
    .Q(net174),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.D(_1551_),
    .Q(net219),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.D(_1552_),
    .Q(net35),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.D(_1553_),
    .Q(net268),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3531_ (.D(_1554_),
    .Q(net143),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.D(_1555_),
    .Q(net244),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3533_ (.D(_1556_),
    .Q(net77),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.D(_1557_),
    .Q(net207),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3535_ (.D(_1558_),
    .Q(net195),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.D(_1560_),
    .Q(net260),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.D(_1561_),
    .Q(net238),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.D(_1562_),
    .Q(net253),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3539_ (.D(_1563_),
    .Q(net129),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.D(_1564_),
    .Q(net18),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.D(_1565_),
    .Q(net185),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3542_ (.D(_1566_),
    .Q(net246),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.D(_1567_),
    .Q(net45),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.D(_1568_),
    .Q(net191),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3545_ (.D(_1569_),
    .Q(net80),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.D(_1571_),
    .Q(net108),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.D(_1572_),
    .Q(net29),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.D(_1573_),
    .Q(net171),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.D(_1574_),
    .Q(net181),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.D(_1575_),
    .Q(net109),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.D(_1576_),
    .Q(net235),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.D(_1577_),
    .Q(net224),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.D(_1578_),
    .Q(net87),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.D(_1579_),
    .Q(net159),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.D(_1580_),
    .Q(net14),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.D(_1582_),
    .Q(net243),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.D(_1583_),
    .Q(net231),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.D(_1584_),
    .Q(net34),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.D(_1585_),
    .Q(net61),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.D(_1586_),
    .Q(net99),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.D(_1587_),
    .Q(net236),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.D(_1588_),
    .Q(net46),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.D(_1589_),
    .Q(net212),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.D(_1590_),
    .Q(net198),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.D(_1591_),
    .Q(net79),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.D(_1593_),
    .Q(net263),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.D(_1594_),
    .Q(net51),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.D(_1595_),
    .Q(net26),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.D(_1596_),
    .Q(net17),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.D(_1597_),
    .Q(net105),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.D(_1598_),
    .Q(net251),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.D(_1599_),
    .Q(net62),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.D(_1600_),
    .Q(net144),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.D(_1601_),
    .Q(net221),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.D(_1602_),
    .Q(net168),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.D(_1604_),
    .Q(net117),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.D(_1605_),
    .Q(net233),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.D(_1606_),
    .Q(net255),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.D(_1607_),
    .Q(net120),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.D(_1608_),
    .Q(net56),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.D(_1609_),
    .Q(net166),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.D(_1610_),
    .Q(net66),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.D(_1611_),
    .Q(net86),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.D(_1612_),
    .Q(net149),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.D(_1613_),
    .Q(net173),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.D(_1360_),
    .Q(net245),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.D(_1361_),
    .Q(net31),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.D(_1362_),
    .Q(net137),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.D(_1363_),
    .Q(net201),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.D(_1364_),
    .Q(net175),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3591_ (.D(_1365_),
    .Q(net42),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.D(_1366_),
    .Q(net202),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.D(_1367_),
    .Q(net122),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3594_ (.D(_1368_),
    .Q(net270),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3595_ (.D(_1369_),
    .Q(net106),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3596_ (.D(_1371_),
    .Q(net49),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3597_ (.D(_1372_),
    .Q(net187),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.D(_1373_),
    .Q(net15),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3599_ (.D(_1374_),
    .Q(net262),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3600_ (.D(_1375_),
    .Q(net192),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.D(_1376_),
    .Q(net38),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3602_ (.D(_1377_),
    .Q(net81),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.D(_1378_),
    .Q(net59),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.D(_1379_),
    .Q(net259),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3605_ (.D(_1380_),
    .Q(net115),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.D(_1382_),
    .Q(net197),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.D(_1383_),
    .Q(net210),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.D(_1384_),
    .Q(net242),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.D(_1385_),
    .Q(net50),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.D(_1386_),
    .Q(net155),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.D(_1387_),
    .Q(net93),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3612_ (.D(_1388_),
    .Q(net158),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3613_ (.D(_1389_),
    .Q(net226),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.D(_1390_),
    .Q(net183),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.D(_1391_),
    .Q(net57),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.D(_1393_),
    .Q(net24),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.D(_1394_),
    .Q(net165),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.D(_1395_),
    .Q(net67),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.D(_1396_),
    .Q(net232),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.D(_1397_),
    .Q(net37),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3621_ (.D(_1398_),
    .Q(net248),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3622_ (.D(_1399_),
    .Q(net134),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3623_ (.D(_1400_),
    .Q(net113),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.D(_1401_),
    .Q(net206),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.D(_1402_),
    .Q(net217),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3626_ (.D(_1404_),
    .Q(net156),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3627_ (.D(_1405_),
    .Q(net214),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3628_ (.D(_1406_),
    .Q(net47),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.D(_1407_),
    .Q(net160),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3630_ (.D(_1408_),
    .Q(net123),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.D(_1409_),
    .Q(net140),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3632_ (.D(_1410_),
    .Q(net127),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.D(_1411_),
    .Q(net131),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.D(_1412_),
    .Q(net228),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.D(_1413_),
    .Q(net145),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.D(_1415_),
    .Q(net220),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.D(_1416_),
    .Q(net40),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.D(_1417_),
    .Q(net199),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.D(_1418_),
    .Q(net265),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.D(_1419_),
    .Q(net148),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.D(_1420_),
    .Q(net204),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.D(_1421_),
    .Q(net167),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.D(_1422_),
    .Q(net114),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.D(_1423_),
    .Q(net142),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.D(_1424_),
    .Q(net196),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.D(_1426_),
    .Q(net75),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.D(_1427_),
    .Q(net73),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.D(_1428_),
    .Q(net126),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.D(_1429_),
    .Q(net118),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.D(_1430_),
    .Q(net111),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.D(_1431_),
    .Q(net256),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.D(_1432_),
    .Q(net19),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.D(_1433_),
    .Q(net194),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.D(_1434_),
    .Q(net128),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.D(_1435_),
    .Q(net176),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.D(_1437_),
    .Q(net213),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.D(_1438_),
    .Q(net239),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.D(_1439_),
    .Q(net247),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.D(_1440_),
    .Q(net250),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3660_ (.D(_1441_),
    .Q(net43),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3661_ (.D(_1442_),
    .Q(net161),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.D(_1443_),
    .Q(net169),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3663_ (.D(_1444_),
    .Q(net227),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3664_ (.D(_1445_),
    .Q(net163),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3665_ (.D(_1446_),
    .Q(net60),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3666_ (.D(_1448_),
    .Q(net179),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3667_ (.D(_1449_),
    .Q(net152),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3668_ (.D(_1450_),
    .Q(net64),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.D(_1451_),
    .Q(net189),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.D(_1452_),
    .Q(net249),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3671_ (.D(_1453_),
    .Q(net90),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.D(_1454_),
    .Q(net178),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3673_ (.D(_1455_),
    .Q(net78),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.D(_1456_),
    .Q(net88),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.D(_1457_),
    .Q(net200),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.D(_1459_),
    .Q(net97),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.D(_1460_),
    .Q(net70),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.D(_1461_),
    .Q(net237),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.D(_1462_),
    .Q(net103),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.D(_1463_),
    .Q(net83),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.D(_1464_),
    .Q(net22),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.D(_1465_),
    .Q(net44),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.D(_1466_),
    .Q(net30),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.D(_1467_),
    .Q(net101),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.D(_1468_),
    .Q(net130),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.D(_1471_),
    .Q(net20),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.D(_1472_),
    .Q(net125),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.D(_1473_),
    .Q(net261),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.D(_1474_),
    .Q(net266),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.D(_1475_),
    .Q(net135),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.D(_1476_),
    .Q(net170),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.D(_1477_),
    .Q(net182),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.D(_1478_),
    .Q(net154),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.D(_1479_),
    .Q(net76),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.D(_1480_),
    .Q(net138),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.D(_1482_),
    .Q(net218),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.D(_1483_),
    .Q(net100),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.D(_1484_),
    .Q(net39),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.D(_1485_),
    .Q(net33),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.D(_1486_),
    .Q(net180),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.D(_1487_),
    .Q(net63),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.D(_1488_),
    .Q(net216),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.D(_1489_),
    .Q(net116),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.D(_1490_),
    .Q(net54),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.D(_1491_),
    .Q(net190),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.D(_1493_),
    .Q(net186),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.D(_1494_),
    .Q(net96),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.D(_1495_),
    .Q(net151),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.D(_1496_),
    .Q(net257),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.D(_1497_),
    .Q(net147),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.D(_1498_),
    .Q(net209),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.D(_1499_),
    .Q(net102),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.D(_1500_),
    .Q(net85),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.D(_1501_),
    .Q(net184),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.D(_1502_),
    .Q(net25),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.D(_1504_),
    .Q(net36),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.D(_1505_),
    .Q(net264),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.D(_1506_),
    .Q(net69),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.D(_1507_),
    .Q(net203),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.D(_1508_),
    .Q(net139),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.D(_1509_),
    .Q(net84),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.D(_1510_),
    .Q(net41),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3723_ (.D(_1511_),
    .Q(net146),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.D(_1512_),
    .Q(net254),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.D(_1513_),
    .Q(net229),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.D(_1515_),
    .Q(net222),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.D(_1516_),
    .Q(net48),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3728_ (.D(_1517_),
    .Q(net52),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3729_ (.D(_1518_),
    .Q(net112),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.D(_1519_),
    .Q(net16),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.D(_1520_),
    .Q(net28),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.D(_1521_),
    .Q(net258),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3733_ (.D(_1522_),
    .Q(net188),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3734_ (.D(_1523_),
    .Q(net164),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3735_ (.D(_1524_),
    .Q(net104),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.D(_1526_),
    .Q(net55),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.D(_1527_),
    .Q(net32),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.D(_1528_),
    .Q(net193),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.D(_1529_),
    .Q(net107),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.D(_1530_),
    .Q(net240),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.D(_1531_),
    .Q(net230),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.D(net4),
    .Q(\input_binary_slice_q[0] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.D(net5),
    .Q(\input_binary_slice_q[1] ),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3744_ (.D(\input_binary_slice_q[0] ),
    .Q(net177),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfxtp_2 _3745_ (.D(\input_binary_slice_q[1] ),
    .Q(net208),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.D(_0515_),
    .Q(\reversed_thermometer[255] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_2 _3747_ (.D(_0001_),
    .Q(\remap_control[0] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_2 _3748_ (.D(_0002_),
    .Q(\remap_control[1] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3749_ (.D(_0000_),
    .Q(\lfsr_q[0] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3750_ (.D(\lfsr_q[0] ),
    .Q(\lfsr_q[1] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3751_ (.D(\lfsr_q[1] ),
    .Q(\lfsr_q[2] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3752_ (.D(\lfsr_q[2] ),
    .Q(\lfsr_q[3] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3753_ (.D(\lfsr_q[3] ),
    .Q(\lfsr_q[4] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3754_ (.D(\lfsr_q[4] ),
    .Q(\lfsr_q[5] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3755_ (.D(\lfsr_q[5] ),
    .Q(\lfsr_q[6] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3756_ (.D(\lfsr_q[6] ),
    .Q(\lfsr_q[7] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3757_ (.D(\lfsr_q[7] ),
    .Q(\lfsr_q[8] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3758_ (.D(\lfsr_q[8] ),
    .Q(\lfsr_q[9] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3759_ (.D(\lfsr_q[9] ),
    .Q(\lfsr_q[10] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3760_ (.D(\lfsr_q[10] ),
    .Q(\lfsr_q[11] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3761_ (.D(\lfsr_q[11] ),
    .Q(\lfsr_q[12] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3762_ (.D(\lfsr_q[12] ),
    .Q(\lfsr_q[13] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 _3763_ (.D(\lfsr_q[13] ),
    .Q(\lfsr_q[14] ),
    .RESET_B(net287),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(rst_ni),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(randomise_en_i),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(en_i),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(input_binary_i[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(input_binary_i[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(input_binary_i[2]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(input_binary_i[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(input_binary_i[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(input_binary_i[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(input_binary_i[6]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(input_binary_i[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(input_binary_i[8]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(input_binary_i[9]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 output14 (.A(net14),
    .X(output_thermometer_o[69]));
 sky130_fd_sc_hd__clkbuf_2 output15 (.A(net15),
    .X(output_thermometer_o[112]));
 sky130_fd_sc_hd__clkbuf_2 output16 (.A(net16),
    .X(output_thermometer_o[244]));
 sky130_fd_sc_hd__clkbuf_2 output17 (.A(net17),
    .X(output_thermometer_o[83]));
 sky130_fd_sc_hd__clkbuf_2 output18 (.A(net18),
    .X(output_thermometer_o[54]));
 sky130_fd_sc_hd__clkbuf_2 output19 (.A(net19),
    .X(output_thermometer_o[166]));
 sky130_fd_sc_hd__clkbuf_2 output20 (.A(net20),
    .X(output_thermometer_o[200]));
 sky130_fd_sc_hd__clkbuf_2 output21 (.A(net21),
    .X(output_thermometer_o[17]));
 sky130_fd_sc_hd__clkbuf_2 output22 (.A(net22),
    .X(output_thermometer_o[195]));
 sky130_fd_sc_hd__clkbuf_2 output23 (.A(net23),
    .X(output_thermometer_o[15]));
 sky130_fd_sc_hd__clkbuf_2 output24 (.A(net24),
    .X(output_thermometer_o[130]));
 sky130_fd_sc_hd__clkbuf_2 output25 (.A(net25),
    .X(output_thermometer_o[229]));
 sky130_fd_sc_hd__clkbuf_2 output26 (.A(net26),
    .X(output_thermometer_o[82]));
 sky130_fd_sc_hd__clkbuf_2 output27 (.A(net27),
    .X(output_thermometer_o[4]));
 sky130_fd_sc_hd__clkbuf_2 output28 (.A(net28),
    .X(output_thermometer_o[245]));
 sky130_fd_sc_hd__clkbuf_2 output29 (.A(net29),
    .X(output_thermometer_o[61]));
 sky130_fd_sc_hd__clkbuf_2 output30 (.A(net30),
    .X(output_thermometer_o[197]));
 sky130_fd_sc_hd__clkbuf_2 output31 (.A(net31),
    .X(output_thermometer_o[101]));
 sky130_fd_sc_hd__clkbuf_2 output32 (.A(net32),
    .X(output_thermometer_o[251]));
 sky130_fd_sc_hd__clkbuf_2 output33 (.A(net33),
    .X(output_thermometer_o[213]));
 sky130_fd_sc_hd__clkbuf_2 output34 (.A(net34),
    .X(output_thermometer_o[72]));
 sky130_fd_sc_hd__clkbuf_2 output35 (.A(net35),
    .X(output_thermometer_o[43]));
 sky130_fd_sc_hd__clkbuf_2 output36 (.A(net36),
    .X(output_thermometer_o[230]));
 sky130_fd_sc_hd__clkbuf_2 output37 (.A(net37),
    .X(output_thermometer_o[134]));
 sky130_fd_sc_hd__clkbuf_2 output38 (.A(net38),
    .X(output_thermometer_o[115]));
 sky130_fd_sc_hd__clkbuf_2 output39 (.A(net39),
    .X(output_thermometer_o[212]));
 sky130_fd_sc_hd__clkbuf_2 output40 (.A(net40),
    .X(output_thermometer_o[151]));
 sky130_fd_sc_hd__clkbuf_2 output41 (.A(net41),
    .X(output_thermometer_o[236]));
 sky130_fd_sc_hd__clkbuf_2 output42 (.A(net42),
    .X(output_thermometer_o[105]));
 sky130_fd_sc_hd__clkbuf_2 output43 (.A(net43),
    .X(output_thermometer_o[174]));
 sky130_fd_sc_hd__clkbuf_2 output44 (.A(net44),
    .X(output_thermometer_o[196]));
 sky130_fd_sc_hd__clkbuf_2 output45 (.A(net45),
    .X(output_thermometer_o[57]));
 sky130_fd_sc_hd__clkbuf_2 output46 (.A(net46),
    .X(output_thermometer_o[76]));
 sky130_fd_sc_hd__clkbuf_2 output47 (.A(net47),
    .X(output_thermometer_o[142]));
 sky130_fd_sc_hd__clkbuf_2 output48 (.A(net48),
    .X(output_thermometer_o[241]));
 sky130_fd_sc_hd__clkbuf_2 output49 (.A(net49),
    .X(output_thermometer_o[110]));
 sky130_fd_sc_hd__clkbuf_2 output50 (.A(net50),
    .X(output_thermometer_o[123]));
 sky130_fd_sc_hd__clkbuf_2 output51 (.A(net51),
    .X(output_thermometer_o[81]));
 sky130_fd_sc_hd__clkbuf_2 output52 (.A(net52),
    .X(output_thermometer_o[242]));
 sky130_fd_sc_hd__clkbuf_2 output53 (.A(net53),
    .X(output_thermometer_o[14]));
 sky130_fd_sc_hd__clkbuf_2 output54 (.A(net54),
    .X(output_thermometer_o[218]));
 sky130_fd_sc_hd__clkbuf_2 output55 (.A(net55),
    .X(output_thermometer_o[250]));
 sky130_fd_sc_hd__clkbuf_2 output56 (.A(net56),
    .X(output_thermometer_o[94]));
 sky130_fd_sc_hd__clkbuf_2 output57 (.A(net57),
    .X(output_thermometer_o[129]));
 sky130_fd_sc_hd__clkbuf_2 output58 (.A(net58),
    .X(output_thermometer_o[9]));
 sky130_fd_sc_hd__clkbuf_2 output59 (.A(net59),
    .X(output_thermometer_o[117]));
 sky130_fd_sc_hd__clkbuf_2 output60 (.A(net60),
    .X(output_thermometer_o[179]));
 sky130_fd_sc_hd__clkbuf_2 output61 (.A(net61),
    .X(output_thermometer_o[73]));
 sky130_fd_sc_hd__clkbuf_2 output62 (.A(net62),
    .X(output_thermometer_o[86]));
 sky130_fd_sc_hd__clkbuf_2 output63 (.A(net63),
    .X(output_thermometer_o[215]));
 sky130_fd_sc_hd__clkbuf_2 output64 (.A(net64),
    .X(output_thermometer_o[182]));
 sky130_fd_sc_hd__clkbuf_2 output65 (.A(net65),
    .X(output_thermometer_o[12]));
 sky130_fd_sc_hd__clkbuf_2 output66 (.A(net66),
    .X(output_thermometer_o[96]));
 sky130_fd_sc_hd__clkbuf_2 output67 (.A(net67),
    .X(output_thermometer_o[132]));
 sky130_fd_sc_hd__clkbuf_2 output68 (.A(net68),
    .X(output_thermometer_o[29]));
 sky130_fd_sc_hd__clkbuf_2 output69 (.A(net69),
    .X(output_thermometer_o[232]));
 sky130_fd_sc_hd__clkbuf_2 output70 (.A(net70),
    .X(output_thermometer_o[191]));
 sky130_fd_sc_hd__clkbuf_2 output71 (.A(net71),
    .X(output_thermometer_o[5]));
 sky130_fd_sc_hd__clkbuf_2 output72 (.A(net72),
    .X(output_thermometer_o[33]));
 sky130_fd_sc_hd__clkbuf_2 output73 (.A(net73),
    .X(output_thermometer_o[161]));
 sky130_fd_sc_hd__clkbuf_2 output74 (.A(net74),
    .X(output_thermometer_o[11]));
 sky130_fd_sc_hd__clkbuf_2 output75 (.A(net75),
    .X(output_thermometer_o[160]));
 sky130_fd_sc_hd__clkbuf_2 output76 (.A(net76),
    .X(output_thermometer_o[208]));
 sky130_fd_sc_hd__clkbuf_2 output77 (.A(net77),
    .X(output_thermometer_o[47]));
 sky130_fd_sc_hd__clkbuf_2 output78 (.A(net78),
    .X(output_thermometer_o[187]));
 sky130_fd_sc_hd__clkbuf_2 output79 (.A(net79),
    .X(output_thermometer_o[79]));
 sky130_fd_sc_hd__clkbuf_2 output80 (.A(net80),
    .X(output_thermometer_o[59]));
 sky130_fd_sc_hd__clkbuf_2 output81 (.A(net81),
    .X(output_thermometer_o[116]));
 sky130_fd_sc_hd__clkbuf_2 output82 (.A(net82),
    .X(output_thermometer_o[30]));
 sky130_fd_sc_hd__clkbuf_2 output83 (.A(net83),
    .X(output_thermometer_o[194]));
 sky130_fd_sc_hd__clkbuf_2 output84 (.A(net84),
    .X(output_thermometer_o[235]));
 sky130_fd_sc_hd__clkbuf_2 output85 (.A(net85),
    .X(output_thermometer_o[227]));
 sky130_fd_sc_hd__clkbuf_2 output86 (.A(net86),
    .X(output_thermometer_o[97]));
 sky130_fd_sc_hd__clkbuf_2 output87 (.A(net87),
    .X(output_thermometer_o[67]));
 sky130_fd_sc_hd__clkbuf_2 output88 (.A(net88),
    .X(output_thermometer_o[188]));
 sky130_fd_sc_hd__clkbuf_2 output89 (.A(net89),
    .X(output_thermometer_o[31]));
 sky130_fd_sc_hd__clkbuf_2 output90 (.A(net90),
    .X(output_thermometer_o[185]));
 sky130_fd_sc_hd__clkbuf_2 output91 (.A(net91),
    .X(output_thermometer_o[20]));
 sky130_fd_sc_hd__clkbuf_2 output92 (.A(net92),
    .X(output_thermometer_o[32]));
 sky130_fd_sc_hd__clkbuf_2 output93 (.A(net93),
    .X(output_thermometer_o[125]));
 sky130_fd_sc_hd__clkbuf_2 output94 (.A(net94),
    .X(output_thermometer_o[7]));
 sky130_fd_sc_hd__clkbuf_2 output95 (.A(net95),
    .X(output_thermometer_o[21]));
 sky130_fd_sc_hd__clkbuf_2 output96 (.A(net96),
    .X(output_thermometer_o[221]));
 sky130_fd_sc_hd__clkbuf_2 output97 (.A(net97),
    .X(output_thermometer_o[190]));
 sky130_fd_sc_hd__clkbuf_2 output98 (.A(net98),
    .X(output_thermometer_o[37]));
 sky130_fd_sc_hd__clkbuf_2 output99 (.A(net99),
    .X(output_thermometer_o[74]));
 sky130_fd_sc_hd__clkbuf_2 output100 (.A(net100),
    .X(output_thermometer_o[211]));
 sky130_fd_sc_hd__clkbuf_2 output101 (.A(net101),
    .X(output_thermometer_o[198]));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(output_thermometer_o[226]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(output_thermometer_o[193]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(output_thermometer_o[249]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(output_thermometer_o[84]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(output_thermometer_o[109]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(output_thermometer_o[253]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(output_thermometer_o[60]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(output_thermometer_o[64]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(output_thermometer_o[23]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(output_thermometer_o[164]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(output_thermometer_o[243]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(output_thermometer_o[137]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(output_thermometer_o[157]));
 sky130_fd_sc_hd__clkbuf_2 output115 (.A(net115),
    .X(output_thermometer_o[119]));
 sky130_fd_sc_hd__clkbuf_2 output116 (.A(net116),
    .X(output_thermometer_o[217]));
 sky130_fd_sc_hd__clkbuf_2 output117 (.A(net117),
    .X(output_thermometer_o[90]));
 sky130_fd_sc_hd__clkbuf_2 output118 (.A(net118),
    .X(output_thermometer_o[163]));
 sky130_fd_sc_hd__clkbuf_2 output119 (.A(net119),
    .X(output_thermometer_o[18]));
 sky130_fd_sc_hd__clkbuf_2 output120 (.A(net120),
    .X(output_thermometer_o[93]));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(output_thermometer_o[26]));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(output_thermometer_o[107]));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(output_thermometer_o[144]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(output_thermometer_o[27]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(output_thermometer_o[201]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(output_thermometer_o[162]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(output_thermometer_o[146]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(output_thermometer_o[168]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(output_thermometer_o[53]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(output_thermometer_o[199]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(output_thermometer_o[147]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(output_thermometer_o[2]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(output_thermometer_o[3]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(output_thermometer_o[136]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(output_thermometer_o[204]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(output_thermometer_o[8]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(output_thermometer_o[102]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(output_thermometer_o[209]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(output_thermometer_o[234]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(output_thermometer_o[145]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(output_thermometer_o[16]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(output_thermometer_o[158]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(output_thermometer_o[45]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(output_thermometer_o[87]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(output_thermometer_o[149]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(output_thermometer_o[237]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(output_thermometer_o[224]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(output_thermometer_o[154]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(output_thermometer_o[98]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(output_thermometer_o[19]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(output_thermometer_o[222]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(output_thermometer_o[181]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(output_thermometer_o[35]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(output_thermometer_o[207]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(output_thermometer_o[124]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(output_thermometer_o[140]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(output_thermometer_o[25]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(output_thermometer_o[126]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(output_thermometer_o[68]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(output_thermometer_o[143]));
 sky130_fd_sc_hd__clkbuf_2 output161 (.A(net161),
    .X(output_thermometer_o[175]));
 sky130_fd_sc_hd__clkbuf_2 output162 (.A(net162),
    .X(output_thermometer_o[13]));
 sky130_fd_sc_hd__clkbuf_2 output163 (.A(net163),
    .X(output_thermometer_o[178]));
 sky130_fd_sc_hd__clkbuf_2 output164 (.A(net164),
    .X(output_thermometer_o[248]));
 sky130_fd_sc_hd__clkbuf_2 output165 (.A(net165),
    .X(output_thermometer_o[131]));
 sky130_fd_sc_hd__clkbuf_2 output166 (.A(net166),
    .X(output_thermometer_o[95]));
 sky130_fd_sc_hd__clkbuf_2 output167 (.A(net167),
    .X(output_thermometer_o[156]));
 sky130_fd_sc_hd__clkbuf_2 output168 (.A(net168),
    .X(output_thermometer_o[89]));
 sky130_fd_sc_hd__clkbuf_2 output169 (.A(net169),
    .X(output_thermometer_o[176]));
 sky130_fd_sc_hd__clkbuf_2 output170 (.A(net170),
    .X(output_thermometer_o[205]));
 sky130_fd_sc_hd__clkbuf_2 output171 (.A(net171),
    .X(output_thermometer_o[62]));
 sky130_fd_sc_hd__clkbuf_2 output172 (.A(net172),
    .X(output_thermometer_o[39]));
 sky130_fd_sc_hd__clkbuf_2 output173 (.A(net173),
    .X(output_thermometer_o[99]));
 sky130_fd_sc_hd__clkbuf_2 output174 (.A(net174),
    .X(output_thermometer_o[41]));
 sky130_fd_sc_hd__clkbuf_2 output175 (.A(net175),
    .X(output_thermometer_o[104]));
 sky130_fd_sc_hd__clkbuf_2 output176 (.A(net176),
    .X(output_thermometer_o[169]));
 sky130_fd_sc_hd__clkbuf_2 output177 (.A(net177),
    .X(output_binary_o[0]));
 sky130_fd_sc_hd__clkbuf_2 output178 (.A(net178),
    .X(output_thermometer_o[186]));
 sky130_fd_sc_hd__clkbuf_2 output179 (.A(net179),
    .X(output_thermometer_o[180]));
 sky130_fd_sc_hd__clkbuf_2 output180 (.A(net180),
    .X(output_thermometer_o[214]));
 sky130_fd_sc_hd__clkbuf_2 output181 (.A(net181),
    .X(output_thermometer_o[63]));
 sky130_fd_sc_hd__clkbuf_2 output182 (.A(net182),
    .X(output_thermometer_o[206]));
 sky130_fd_sc_hd__clkbuf_2 output183 (.A(net183),
    .X(output_thermometer_o[128]));
 sky130_fd_sc_hd__clkbuf_2 output184 (.A(net184),
    .X(output_thermometer_o[228]));
 sky130_fd_sc_hd__clkbuf_2 output185 (.A(net185),
    .X(output_thermometer_o[55]));
 sky130_fd_sc_hd__clkbuf_2 output186 (.A(net186),
    .X(output_thermometer_o[220]));
 sky130_fd_sc_hd__clkbuf_2 output187 (.A(net187),
    .X(output_thermometer_o[111]));
 sky130_fd_sc_hd__clkbuf_2 output188 (.A(net188),
    .X(output_thermometer_o[247]));
 sky130_fd_sc_hd__clkbuf_2 output189 (.A(net189),
    .X(output_thermometer_o[183]));
 sky130_fd_sc_hd__clkbuf_2 output190 (.A(net190),
    .X(output_thermometer_o[219]));
 sky130_fd_sc_hd__clkbuf_2 output191 (.A(net191),
    .X(output_thermometer_o[58]));
 sky130_fd_sc_hd__clkbuf_2 output192 (.A(net192),
    .X(output_thermometer_o[114]));
 sky130_fd_sc_hd__clkbuf_2 output193 (.A(net193),
    .X(output_thermometer_o[252]));
 sky130_fd_sc_hd__clkbuf_2 output194 (.A(net194),
    .X(output_thermometer_o[167]));
 sky130_fd_sc_hd__clkbuf_2 output195 (.A(net195),
    .X(output_thermometer_o[49]));
 sky130_fd_sc_hd__clkbuf_2 output196 (.A(net196),
    .X(output_thermometer_o[159]));
 sky130_fd_sc_hd__clkbuf_2 output197 (.A(net197),
    .X(output_thermometer_o[120]));
 sky130_fd_sc_hd__clkbuf_2 output198 (.A(net198),
    .X(output_thermometer_o[78]));
 sky130_fd_sc_hd__clkbuf_2 output199 (.A(net199),
    .X(output_thermometer_o[152]));
 sky130_fd_sc_hd__clkbuf_2 output200 (.A(net200),
    .X(output_thermometer_o[189]));
 sky130_fd_sc_hd__clkbuf_2 output201 (.A(net201),
    .X(output_thermometer_o[103]));
 sky130_fd_sc_hd__clkbuf_2 output202 (.A(net202),
    .X(output_thermometer_o[106]));
 sky130_fd_sc_hd__clkbuf_2 output203 (.A(net203),
    .X(output_thermometer_o[233]));
 sky130_fd_sc_hd__clkbuf_2 output204 (.A(net204),
    .X(output_thermometer_o[155]));
 sky130_fd_sc_hd__clkbuf_2 output205 (.A(net205),
    .X(output_thermometer_o[34]));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(output_thermometer_o[138]));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(output_thermometer_o[48]));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(output_binary_o[1]));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(output_thermometer_o[225]));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(output_thermometer_o[121]));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(output_thermometer_o[10]));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(output_thermometer_o[77]));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(output_thermometer_o[170]));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(output_thermometer_o[141]));
 sky130_fd_sc_hd__clkbuf_2 output215 (.A(net215),
    .X(output_thermometer_o[40]));
 sky130_fd_sc_hd__clkbuf_2 output216 (.A(net216),
    .X(output_thermometer_o[216]));
 sky130_fd_sc_hd__clkbuf_2 output217 (.A(net217),
    .X(output_thermometer_o[139]));
 sky130_fd_sc_hd__clkbuf_2 output218 (.A(net218),
    .X(output_thermometer_o[210]));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(output_thermometer_o[42]));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(output_thermometer_o[150]));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(output_thermometer_o[88]));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net222),
    .X(output_thermometer_o[240]));
 sky130_fd_sc_hd__clkbuf_2 output223 (.A(net223),
    .X(output_thermometer_o[1]));
 sky130_fd_sc_hd__clkbuf_2 output224 (.A(net224),
    .X(output_thermometer_o[66]));
 sky130_fd_sc_hd__clkbuf_2 output225 (.A(net225),
    .X(output_thermometer_o[36]));
 sky130_fd_sc_hd__clkbuf_2 output226 (.A(net226),
    .X(output_thermometer_o[127]));
 sky130_fd_sc_hd__clkbuf_2 output227 (.A(net227),
    .X(output_thermometer_o[177]));
 sky130_fd_sc_hd__clkbuf_2 output228 (.A(net228),
    .X(output_thermometer_o[148]));
 sky130_fd_sc_hd__clkbuf_2 output229 (.A(net229),
    .X(output_thermometer_o[239]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(output_thermometer_o[255]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(output_thermometer_o[71]));
 sky130_fd_sc_hd__clkbuf_2 output232 (.A(net232),
    .X(output_thermometer_o[133]));
 sky130_fd_sc_hd__clkbuf_2 output233 (.A(net233),
    .X(output_thermometer_o[91]));
 sky130_fd_sc_hd__clkbuf_2 output234 (.A(net234),
    .X(output_thermometer_o[22]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net235),
    .X(output_thermometer_o[65]));
 sky130_fd_sc_hd__clkbuf_2 output236 (.A(net236),
    .X(output_thermometer_o[75]));
 sky130_fd_sc_hd__clkbuf_2 output237 (.A(net237),
    .X(output_thermometer_o[192]));
 sky130_fd_sc_hd__clkbuf_2 output238 (.A(net238),
    .X(output_thermometer_o[51]));
 sky130_fd_sc_hd__clkbuf_2 output239 (.A(net239),
    .X(output_thermometer_o[171]));
 sky130_fd_sc_hd__clkbuf_2 output240 (.A(net240),
    .X(output_thermometer_o[254]));
 sky130_fd_sc_hd__clkbuf_2 output241 (.A(net241),
    .X(output_thermometer_o[28]));
 sky130_fd_sc_hd__clkbuf_2 output242 (.A(net242),
    .X(output_thermometer_o[122]));
 sky130_fd_sc_hd__clkbuf_2 output243 (.A(net243),
    .X(output_thermometer_o[70]));
 sky130_fd_sc_hd__clkbuf_2 output244 (.A(net244),
    .X(output_thermometer_o[46]));
 sky130_fd_sc_hd__clkbuf_2 output245 (.A(net245),
    .X(output_thermometer_o[100]));
 sky130_fd_sc_hd__clkbuf_2 output246 (.A(net246),
    .X(output_thermometer_o[56]));
 sky130_fd_sc_hd__clkbuf_2 output247 (.A(net247),
    .X(output_thermometer_o[172]));
 sky130_fd_sc_hd__clkbuf_2 output248 (.A(net248),
    .X(output_thermometer_o[135]));
 sky130_fd_sc_hd__clkbuf_2 output249 (.A(net249),
    .X(output_thermometer_o[184]));
 sky130_fd_sc_hd__clkbuf_2 output250 (.A(net250),
    .X(output_thermometer_o[173]));
 sky130_fd_sc_hd__clkbuf_2 output251 (.A(net251),
    .X(output_thermometer_o[85]));
 sky130_fd_sc_hd__clkbuf_2 output252 (.A(net252),
    .X(output_thermometer_o[38]));
 sky130_fd_sc_hd__clkbuf_2 output253 (.A(net253),
    .X(output_thermometer_o[52]));
 sky130_fd_sc_hd__clkbuf_2 output254 (.A(net254),
    .X(output_thermometer_o[238]));
 sky130_fd_sc_hd__clkbuf_2 output255 (.A(net255),
    .X(output_thermometer_o[92]));
 sky130_fd_sc_hd__clkbuf_2 output256 (.A(net256),
    .X(output_thermometer_o[165]));
 sky130_fd_sc_hd__clkbuf_2 output257 (.A(net257),
    .X(output_thermometer_o[223]));
 sky130_fd_sc_hd__clkbuf_2 output258 (.A(net258),
    .X(output_thermometer_o[246]));
 sky130_fd_sc_hd__clkbuf_2 output259 (.A(net259),
    .X(output_thermometer_o[118]));
 sky130_fd_sc_hd__clkbuf_2 output260 (.A(net260),
    .X(output_thermometer_o[50]));
 sky130_fd_sc_hd__clkbuf_2 output261 (.A(net261),
    .X(output_thermometer_o[202]));
 sky130_fd_sc_hd__clkbuf_2 output262 (.A(net262),
    .X(output_thermometer_o[113]));
 sky130_fd_sc_hd__clkbuf_2 output263 (.A(net263),
    .X(output_thermometer_o[80]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(output_thermometer_o[231]));
 sky130_fd_sc_hd__clkbuf_2 output265 (.A(net265),
    .X(output_thermometer_o[153]));
 sky130_fd_sc_hd__clkbuf_2 output266 (.A(net266),
    .X(output_thermometer_o[203]));
 sky130_fd_sc_hd__clkbuf_2 output267 (.A(net267),
    .X(output_thermometer_o[6]));
 sky130_fd_sc_hd__clkbuf_2 output268 (.A(net268),
    .X(output_thermometer_o[44]));
 sky130_fd_sc_hd__clkbuf_2 output269 (.A(net269),
    .X(output_thermometer_o[0]));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(output_thermometer_o[108]));
 sky130_fd_sc_hd__clkbuf_2 output271 (.A(net271),
    .X(output_thermometer_o[24]));
 sky130_fd_sc_hd__clkbuf_2 output272 (.A(net272),
    .X(en_o));
 sky130_fd_sc_hd__buf_8 repeater273 (.A(net286),
    .X(net273));
 sky130_fd_sc_hd__buf_6 repeater274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_8 repeater275 (.A(net277),
    .X(net275));
 sky130_fd_sc_hd__buf_8 repeater276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_8 repeater277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_8 repeater278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_8 repeater279 (.A(net281),
    .X(net279));
 sky130_fd_sc_hd__buf_8 repeater280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_8 repeater281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_6 repeater282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__buf_6 repeater283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_6 repeater284 (.A(net286),
    .X(net284));
 sky130_fd_sc_hd__buf_8 repeater285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_8 repeater286 (.A(_0227_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_clk_i (.A(clknet_1_0_0_clk_i),
    .X(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_clk_i (.A(clknet_1_0_0_clk_i),
    .X(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_clk_i (.A(clknet_1_1_0_clk_i),
    .X(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_clk_i (.A(clknet_1_1_0_clk_i),
    .X(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net1),
    .X(net287));
endmodule
