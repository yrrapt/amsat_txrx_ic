* Generic MOS noise characterisation netlist

.param temp=27
.temp 27

* .lib "sky130_fd_pr/models/sky130.lib.spice" tt
.include "sky130_fd_pr/models/corners/tt.spice"

.param id=10u
.param vds=1.8
.param vdd=1.8
.param vbs=0
.param l=0.15
.param vctl=-10

* XMcurr net1 gate vdd vdd sky130_fd_pr__pfet_01v8_lvt w=1 l=1 m=1



XM vd vg 0 vb sky130_fd_pr__nfet_01v8_lvt w=1 l=1 m=1

Bgs vg 0 V=min(i(Vds)*1e9,vdd)
BId 0 vd I=10**v(vctl)
Vds vd_ 0 DC={vds} AC=0
Vbs vb 0 {vbs}
Vctl vctl 0 {vctl}

Vdmeas vd vd_
Hccvs out 0 Vdmeas 1

* Vdd vdd 0 {vdd} 
* Vgate vdd gate DC=0.8 AC=1
* Vout net1 0 0.7

* specify op paramters to save
.save all @m.xm.msky130_fd_pr__nfet_01v8_lvt[vdsat] @m.xm.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm.msky130_fd_pr__nfet_01v8_lvt[gm] @m.xm.msky130_fd_pr__nfet_01v8_lvt[id]


* specify the simulations
* .dc Vctl -10 -3 0.01
* .dc Vctl -10 -3 0.01

.op
.noise v(out) Vds dec 10 1 100000Meg

.control
  run
  setplot op1
  write spiceinterface_temp_dc1.raw
  setplot noise1
  write spiceinterface_temp_noise1.raw
  * quit
.endc


* .control
* let start_vctl = -10
* let stop_vctl = -3
* let delta_vctl = 0.01
* let act_vctl = start_vctl

* while act_vctl le stop_vctl
    
*     * start a new simulation
*     alter vctl act_vctl
*     run

*     * save the results
*     setplot dc1
*     write spiceinterface_temp_dc.raw
*     setplot noise1
*     write spiceinterface_temp_noise.raw
*     set appendwrite

*     * move to next step
*     let act_vctl = act_vctl + delta_vctl
* end
* .endc


.end