VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dac_digital_interface
  CLASS BLOCK ;
  FOREIGN dac_digital_interface ;
  ORIGIN 0.000 0.000 ;
  SIZE 270.000 BY 210.000 ;
  PIN output_thermometer_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.570 208.350 5.710 210.000 ;
    END
  END output_thermometer_o[69]
  PIN output_thermometer_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.570 0.000 5.710 1.090 ;
    END
  END output_thermometer_o[112]
  PIN output_thermometer_o[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.950 208.350 7.090 210.000 ;
    END
  END output_thermometer_o[244]
  PIN output_thermometer_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.950 0.000 7.090 1.090 ;
    END
  END output_thermometer_o[83]
  PIN output_thermometer_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.330 208.350 8.470 210.000 ;
    END
  END output_thermometer_o[54]
  PIN output_thermometer_o[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.330 0.000 8.470 1.090 ;
    END
  END output_thermometer_o[166]
  PIN output_thermometer_o[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.710 208.350 9.850 210.000 ;
    END
  END output_thermometer_o[200]
  PIN output_thermometer_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.710 0.000 9.850 1.090 ;
    END
  END output_thermometer_o[17]
  PIN output_thermometer_o[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.090 208.350 11.230 210.000 ;
    END
  END output_thermometer_o[195]
  PIN output_thermometer_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.090 0.000 11.230 1.090 ;
    END
  END output_thermometer_o[15]
  PIN output_thermometer_o[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.470 208.350 12.610 210.000 ;
    END
  END output_thermometer_o[130]
  PIN output_thermometer_o[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.470 0.000 12.610 0.410 ;
    END
  END output_thermometer_o[229]
  PIN output_thermometer_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.850 208.350 13.990 210.000 ;
    END
  END output_thermometer_o[82]
  PIN output_thermometer_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.850 0.000 13.990 1.090 ;
    END
  END output_thermometer_o[4]
  PIN output_thermometer_o[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.230 208.350 15.370 210.000 ;
    END
  END output_thermometer_o[245]
  PIN output_thermometer_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.230 0.000 15.370 1.090 ;
    END
  END output_thermometer_o[61]
  PIN output_thermometer_o[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.610 208.350 16.750 210.000 ;
    END
  END output_thermometer_o[197]
  PIN output_thermometer_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.610 0.000 16.750 1.090 ;
    END
  END output_thermometer_o[101]
  PIN output_thermometer_o[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.990 208.350 18.130 210.000 ;
    END
  END output_thermometer_o[251]
  PIN output_thermometer_o[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.990 0.000 18.130 1.090 ;
    END
  END output_thermometer_o[213]
  PIN output_thermometer_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.370 208.350 19.510 210.000 ;
    END
  END output_thermometer_o[72]
  PIN output_thermometer_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.370 0.000 19.510 0.410 ;
    END
  END output_thermometer_o[43]
  PIN output_thermometer_o[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.750 208.720 20.890 210.000 ;
    END
  END output_thermometer_o[230]
  PIN output_thermometer_o[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.750 0.000 20.890 0.410 ;
    END
  END output_thermometer_o[134]
  PIN output_thermometer_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.130 209.060 22.270 210.000 ;
    END
  END output_thermometer_o[115]
  PIN output_thermometer_o[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.130 0.000 22.270 0.410 ;
    END
  END output_thermometer_o[212]
  PIN output_thermometer_o[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.510 208.350 23.650 210.000 ;
    END
  END output_thermometer_o[151]
  PIN output_thermometer_o[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.510 0.000 23.650 0.410 ;
    END
  END output_thermometer_o[236]
  PIN output_thermometer_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.890 208.350 25.030 210.000 ;
    END
  END output_thermometer_o[105]
  PIN output_thermometer_o[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.890 0.000 25.030 0.410 ;
    END
  END output_thermometer_o[174]
  PIN output_thermometer_o[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.270 208.350 26.410 210.000 ;
    END
  END output_thermometer_o[196]
  PIN output_thermometer_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.270 0.000 26.410 1.090 ;
    END
  END output_thermometer_o[57]
  PIN output_thermometer_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.650 208.350 27.790 210.000 ;
    END
  END output_thermometer_o[76]
  PIN output_thermometer_o[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.650 0.000 27.790 1.060 ;
    END
  END output_thermometer_o[142]
  PIN output_thermometer_o[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.030 208.350 29.170 210.000 ;
    END
  END output_thermometer_o[241]
  PIN output_thermometer_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.030 0.000 29.170 1.090 ;
    END
  END output_thermometer_o[110]
  PIN output_thermometer_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.410 208.350 30.550 210.000 ;
    END
  END output_thermometer_o[123]
  PIN output_thermometer_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.410 0.000 30.550 0.410 ;
    END
  END output_thermometer_o[81]
  PIN output_thermometer_o[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.790 208.350 31.930 210.000 ;
    END
  END output_thermometer_o[242]
  PIN output_thermometer_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.790 0.000 31.930 1.060 ;
    END
  END output_thermometer_o[14]
  PIN output_thermometer_o[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.170 208.350 33.310 210.000 ;
    END
  END output_thermometer_o[218]
  PIN output_thermometer_o[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.170 0.000 33.310 1.090 ;
    END
  END output_thermometer_o[250]
  PIN output_thermometer_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.550 208.350 34.690 210.000 ;
    END
  END output_thermometer_o[94]
  PIN output_thermometer_o[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.550 0.000 34.690 0.410 ;
    END
  END output_thermometer_o[129]
  PIN output_thermometer_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.930 208.350 36.070 210.000 ;
    END
  END output_thermometer_o[9]
  PIN output_thermometer_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.930 0.000 36.070 0.410 ;
    END
  END output_thermometer_o[117]
  PIN output_thermometer_o[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.310 208.350 37.450 210.000 ;
    END
  END output_thermometer_o[179]
  PIN output_thermometer_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.310 0.000 37.450 0.410 ;
    END
  END output_thermometer_o[73]
  PIN output_thermometer_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.690 208.350 38.830 210.000 ;
    END
  END output_thermometer_o[86]
  PIN output_thermometer_o[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.690 0.000 38.830 1.090 ;
    END
  END output_thermometer_o[215]
  PIN output_thermometer_o[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.070 208.350 40.210 210.000 ;
    END
  END output_thermometer_o[182]
  PIN output_thermometer_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.070 0.000 40.210 1.090 ;
    END
  END output_thermometer_o[12]
  PIN output_thermometer_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.450 208.350 41.590 210.000 ;
    END
  END output_thermometer_o[96]
  PIN output_thermometer_o[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.450 0.000 41.590 0.410 ;
    END
  END output_thermometer_o[132]
  PIN output_thermometer_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.830 208.350 42.970 210.000 ;
    END
  END output_thermometer_o[29]
  PIN output_thermometer_o[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.830 0.000 42.970 0.410 ;
    END
  END output_thermometer_o[232]
  PIN output_thermometer_o[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.210 208.350 44.350 210.000 ;
    END
  END output_thermometer_o[191]
  PIN output_thermometer_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.210 0.000 44.350 0.410 ;
    END
  END output_thermometer_o[5]
  PIN output_thermometer_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.590 208.350 45.730 210.000 ;
    END
  END output_thermometer_o[33]
  PIN output_thermometer_o[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.590 0.000 45.730 0.410 ;
    END
  END output_thermometer_o[161]
  PIN output_thermometer_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.970 208.350 47.110 210.000 ;
    END
  END output_thermometer_o[11]
  PIN output_thermometer_o[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.970 0.000 47.110 1.090 ;
    END
  END output_thermometer_o[160]
  PIN output_thermometer_o[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.350 208.350 48.490 210.000 ;
    END
  END output_thermometer_o[208]
  PIN output_thermometer_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.350 0.000 48.490 0.410 ;
    END
  END output_thermometer_o[47]
  PIN output_thermometer_o[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.730 208.350 49.870 210.000 ;
    END
  END output_thermometer_o[187]
  PIN output_thermometer_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.730 0.000 49.870 0.410 ;
    END
  END output_thermometer_o[79]
  PIN output_thermometer_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.110 208.350 51.250 210.000 ;
    END
  END output_thermometer_o[59]
  PIN output_thermometer_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.110 0.000 51.250 0.410 ;
    END
  END output_thermometer_o[116]
  PIN output_thermometer_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.490 209.030 52.630 210.000 ;
    END
  END output_thermometer_o[30]
  PIN output_thermometer_o[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.490 0.000 52.630 0.410 ;
    END
  END output_thermometer_o[194]
  PIN output_thermometer_o[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.870 208.350 54.010 210.000 ;
    END
  END output_thermometer_o[235]
  PIN output_thermometer_o[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.870 0.000 54.010 0.410 ;
    END
  END output_thermometer_o[227]
  PIN output_thermometer_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.250 208.350 55.390 210.000 ;
    END
  END output_thermometer_o[97]
  PIN output_thermometer_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.250 0.000 55.390 1.090 ;
    END
  END output_thermometer_o[67]
  PIN output_thermometer_o[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.630 208.350 56.770 210.000 ;
    END
  END output_thermometer_o[188]
  PIN output_thermometer_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.630 0.000 56.770 0.410 ;
    END
  END output_thermometer_o[31]
  PIN output_thermometer_o[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.010 208.350 58.150 210.000 ;
    END
  END output_thermometer_o[185]
  PIN output_thermometer_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.010 0.000 58.150 0.410 ;
    END
  END output_thermometer_o[20]
  PIN output_thermometer_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.390 208.350 59.530 210.000 ;
    END
  END output_thermometer_o[32]
  PIN output_thermometer_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.390 0.000 59.530 1.090 ;
    END
  END output_thermometer_o[125]
  PIN output_thermometer_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.770 208.350 60.910 210.000 ;
    END
  END output_thermometer_o[7]
  PIN output_thermometer_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.770 0.000 60.910 0.410 ;
    END
  END output_thermometer_o[21]
  PIN output_thermometer_o[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.150 208.350 62.290 210.000 ;
    END
  END output_thermometer_o[221]
  PIN output_thermometer_o[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.150 0.000 62.290 0.720 ;
    END
  END output_thermometer_o[190]
  PIN output_thermometer_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.530 208.350 63.670 210.000 ;
    END
  END output_thermometer_o[37]
  PIN output_thermometer_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.530 0.000 63.670 1.060 ;
    END
  END output_thermometer_o[74]
  PIN output_thermometer_o[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.910 208.350 65.050 210.000 ;
    END
  END output_thermometer_o[211]
  PIN output_thermometer_o[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.910 0.000 65.050 0.410 ;
    END
  END output_thermometer_o[198]
  PIN output_thermometer_o[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.290 208.350 66.430 210.000 ;
    END
  END output_thermometer_o[226]
  PIN output_thermometer_o[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.290 0.000 66.430 1.090 ;
    END
  END output_thermometer_o[193]
  PIN output_thermometer_o[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.670 208.350 67.810 210.000 ;
    END
  END output_thermometer_o[249]
  PIN output_thermometer_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.670 0.000 67.810 1.090 ;
    END
  END output_thermometer_o[84]
  PIN output_thermometer_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.050 208.350 69.190 210.000 ;
    END
  END output_thermometer_o[109]
  PIN output_thermometer_o[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.050 0.000 69.190 1.090 ;
    END
  END output_thermometer_o[253]
  PIN output_thermometer_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.430 208.350 70.570 210.000 ;
    END
  END output_thermometer_o[60]
  PIN output_thermometer_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.430 0.000 70.570 1.090 ;
    END
  END output_thermometer_o[64]
  PIN output_thermometer_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.810 208.350 71.950 210.000 ;
    END
  END output_thermometer_o[23]
  PIN output_thermometer_o[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.810 0.000 71.950 1.090 ;
    END
  END output_thermometer_o[164]
  PIN output_thermometer_o[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.190 208.350 73.330 210.000 ;
    END
  END output_thermometer_o[243]
  PIN output_thermometer_o[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.190 0.000 73.330 0.410 ;
    END
  END output_thermometer_o[137]
  PIN output_thermometer_o[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.570 208.350 74.710 210.000 ;
    END
  END output_thermometer_o[157]
  PIN output_thermometer_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.570 0.000 74.710 0.410 ;
    END
  END output_thermometer_o[119]
  PIN output_thermometer_o[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.950 208.350 76.090 210.000 ;
    END
  END output_thermometer_o[217]
  PIN output_thermometer_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.950 0.000 76.090 0.410 ;
    END
  END output_thermometer_o[90]
  PIN output_thermometer_o[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.330 208.350 77.470 210.000 ;
    END
  END output_thermometer_o[163]
  PIN output_thermometer_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.330 0.000 77.470 0.410 ;
    END
  END output_thermometer_o[18]
  PIN output_thermometer_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.710 208.350 78.850 210.000 ;
    END
  END output_thermometer_o[93]
  PIN output_thermometer_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.710 0.000 78.850 1.260 ;
    END
  END output_thermometer_o[26]
  PIN output_thermometer_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.090 208.350 80.230 210.000 ;
    END
  END output_thermometer_o[107]
  PIN output_thermometer_o[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.090 0.000 80.230 1.090 ;
    END
  END output_thermometer_o[144]
  PIN output_thermometer_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.470 208.350 81.610 210.000 ;
    END
  END output_thermometer_o[27]
  PIN output_thermometer_o[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.470 0.000 81.610 1.090 ;
    END
  END output_thermometer_o[201]
  PIN output_thermometer_o[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.850 208.350 82.990 210.000 ;
    END
  END output_thermometer_o[162]
  PIN output_thermometer_o[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.850 0.000 82.990 0.410 ;
    END
  END output_thermometer_o[146]
  PIN output_thermometer_o[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.230 208.350 84.370 210.000 ;
    END
  END output_thermometer_o[168]
  PIN output_thermometer_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.230 0.000 84.370 0.410 ;
    END
  END output_thermometer_o[53]
  PIN output_thermometer_o[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.610 208.350 85.750 210.000 ;
    END
  END output_thermometer_o[199]
  PIN output_thermometer_o[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.610 0.000 85.750 1.090 ;
    END
  END output_thermometer_o[147]
  PIN output_thermometer_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.990 209.030 87.130 210.000 ;
    END
  END output_thermometer_o[2]
  PIN output_thermometer_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.990 0.000 87.130 1.090 ;
    END
  END output_thermometer_o[3]
  PIN output_thermometer_o[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.370 208.350 88.510 210.000 ;
    END
  END output_thermometer_o[136]
  PIN output_thermometer_o[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.370 0.000 88.510 1.090 ;
    END
  END output_thermometer_o[204]
  PIN output_thermometer_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.750 208.350 89.890 210.000 ;
    END
  END output_thermometer_o[8]
  PIN output_thermometer_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.750 0.000 89.890 1.090 ;
    END
  END output_thermometer_o[102]
  PIN output_thermometer_o[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.130 208.350 91.270 210.000 ;
    END
  END output_thermometer_o[209]
  PIN output_thermometer_o[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.130 0.000 91.270 1.090 ;
    END
  END output_thermometer_o[234]
  PIN output_thermometer_o[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.510 208.350 92.650 210.000 ;
    END
  END output_thermometer_o[145]
  PIN output_thermometer_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.510 0.000 92.650 0.410 ;
    END
  END output_thermometer_o[16]
  PIN output_thermometer_o[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.890 208.350 94.030 210.000 ;
    END
  END output_thermometer_o[158]
  PIN output_thermometer_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.890 0.000 94.030 0.410 ;
    END
  END output_thermometer_o[45]
  PIN output_thermometer_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.270 208.350 95.410 210.000 ;
    END
  END output_thermometer_o[87]
  PIN output_thermometer_o[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.270 0.000 95.410 1.090 ;
    END
  END output_thermometer_o[149]
  PIN output_thermometer_o[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.650 209.060 96.790 210.000 ;
    END
  END output_thermometer_o[237]
  PIN output_thermometer_o[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.650 0.000 96.790 0.410 ;
    END
  END output_thermometer_o[224]
  PIN output_thermometer_o[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.030 208.720 98.170 210.000 ;
    END
  END output_thermometer_o[154]
  PIN output_thermometer_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.030 0.000 98.170 1.260 ;
    END
  END output_thermometer_o[98]
  PIN output_thermometer_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.410 208.350 99.550 210.000 ;
    END
  END output_thermometer_o[19]
  PIN output_thermometer_o[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.410 0.000 99.550 0.410 ;
    END
  END output_thermometer_o[222]
  PIN output_thermometer_o[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.790 208.350 100.930 210.000 ;
    END
  END output_thermometer_o[181]
  PIN output_thermometer_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.790 0.000 100.930 0.410 ;
    END
  END output_thermometer_o[35]
  PIN output_thermometer_o[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.170 208.350 102.310 210.000 ;
    END
  END output_thermometer_o[207]
  PIN output_thermometer_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.170 0.000 102.310 0.410 ;
    END
  END output_thermometer_o[124]
  PIN output_thermometer_o[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.550 208.350 103.690 210.000 ;
    END
  END output_thermometer_o[140]
  PIN output_thermometer_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.550 0.000 103.690 0.410 ;
    END
  END output_thermometer_o[25]
  PIN output_thermometer_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.930 208.350 105.070 210.000 ;
    END
  END output_thermometer_o[126]
  PIN output_thermometer_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.930 0.000 105.070 1.090 ;
    END
  END output_thermometer_o[68]
  PIN output_thermometer_o[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.310 208.350 106.450 210.000 ;
    END
  END output_thermometer_o[143]
  PIN output_thermometer_o[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.310 0.000 106.450 1.260 ;
    END
  END output_thermometer_o[175]
  PIN output_thermometer_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.690 208.350 107.830 210.000 ;
    END
  END output_thermometer_o[13]
  PIN output_thermometer_o[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.690 0.000 107.830 1.090 ;
    END
  END output_thermometer_o[178]
  PIN output_thermometer_o[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.070 208.350 109.210 210.000 ;
    END
  END output_thermometer_o[248]
  PIN output_thermometer_o[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.070 0.000 109.210 0.410 ;
    END
  END output_thermometer_o[131]
  PIN output_thermometer_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.450 208.720 110.590 210.000 ;
    END
  END output_thermometer_o[95]
  PIN output_thermometer_o[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.450 0.000 110.590 0.410 ;
    END
  END output_thermometer_o[156]
  PIN output_thermometer_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.830 208.350 111.970 210.000 ;
    END
  END output_thermometer_o[89]
  PIN output_thermometer_o[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.830 0.000 111.970 1.090 ;
    END
  END output_thermometer_o[176]
  PIN output_thermometer_o[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.210 208.350 113.350 210.000 ;
    END
  END output_thermometer_o[205]
  PIN output_thermometer_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.210 0.000 113.350 1.090 ;
    END
  END output_thermometer_o[62]
  PIN output_thermometer_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.590 208.350 114.730 210.000 ;
    END
  END output_thermometer_o[39]
  PIN output_thermometer_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.590 0.000 114.730 1.260 ;
    END
  END output_thermometer_o[99]
  PIN output_thermometer_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.970 208.350 116.110 210.000 ;
    END
  END output_thermometer_o[41]
  PIN output_thermometer_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.970 0.000 116.110 1.060 ;
    END
  END output_thermometer_o[104]
  PIN output_thermometer_o[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.350 208.350 117.490 210.000 ;
    END
  END output_thermometer_o[169]
  PIN output_binary_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.350 0.000 117.490 0.410 ;
    END
  END output_binary_o[0]
  PIN output_thermometer_o[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.730 208.350 118.870 210.000 ;
    END
  END output_thermometer_o[186]
  PIN output_thermometer_o[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.730 0.000 118.870 0.410 ;
    END
  END output_thermometer_o[180]
  PIN output_thermometer_o[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.110 208.350 120.250 210.000 ;
    END
  END output_thermometer_o[214]
  PIN output_thermometer_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.110 0.000 120.250 0.410 ;
    END
  END output_thermometer_o[63]
  PIN output_thermometer_o[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.490 208.350 121.630 210.000 ;
    END
  END output_thermometer_o[206]
  PIN output_thermometer_o[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.490 0.000 121.630 1.090 ;
    END
  END output_thermometer_o[128]
  PIN output_thermometer_o[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.870 208.350 123.010 210.000 ;
    END
  END output_thermometer_o[228]
  PIN output_thermometer_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.870 0.000 123.010 0.410 ;
    END
  END output_thermometer_o[55]
  PIN output_thermometer_o[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.250 208.350 124.390 210.000 ;
    END
  END output_thermometer_o[220]
  PIN output_thermometer_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.250 0.000 124.390 1.090 ;
    END
  END output_thermometer_o[111]
  PIN output_thermometer_o[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.630 208.350 125.770 210.000 ;
    END
  END output_thermometer_o[247]
  PIN output_thermometer_o[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.630 0.000 125.770 1.090 ;
    END
  END output_thermometer_o[183]
  PIN output_thermometer_o[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.010 208.350 127.150 210.000 ;
    END
  END output_thermometer_o[219]
  PIN output_thermometer_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.010 0.000 127.150 0.410 ;
    END
  END output_thermometer_o[58]
  PIN output_thermometer_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.390 208.350 128.530 210.000 ;
    END
  END output_thermometer_o[114]
  PIN output_thermometer_o[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.390 0.000 128.530 0.720 ;
    END
  END output_thermometer_o[252]
  PIN output_thermometer_o[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.770 208.350 129.910 210.000 ;
    END
  END output_thermometer_o[167]
  PIN output_thermometer_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.770 0.000 129.910 1.090 ;
    END
  END output_thermometer_o[49]
  PIN output_thermometer_o[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.150 208.350 131.290 210.000 ;
    END
  END output_thermometer_o[159]
  PIN output_thermometer_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.150 0.000 131.290 0.410 ;
    END
  END output_thermometer_o[120]
  PIN output_thermometer_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.530 208.720 132.670 210.000 ;
    END
  END output_thermometer_o[78]
  PIN output_thermometer_o[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.530 0.000 132.670 1.090 ;
    END
  END output_thermometer_o[152]
  PIN output_thermometer_o[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.910 208.350 134.050 210.000 ;
    END
  END output_thermometer_o[189]
  PIN output_thermometer_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.910 0.000 134.050 1.090 ;
    END
  END output_thermometer_o[103]
  PIN output_thermometer_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.290 208.350 135.430 210.000 ;
    END
  END output_thermometer_o[106]
  PIN output_thermometer_o[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.290 0.000 135.430 0.410 ;
    END
  END output_thermometer_o[233]
  PIN output_thermometer_o[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.670 208.350 136.810 210.000 ;
    END
  END output_thermometer_o[155]
  PIN output_thermometer_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.670 0.000 136.810 0.410 ;
    END
  END output_thermometer_o[34]
  PIN output_thermometer_o[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.050 208.350 138.190 210.000 ;
    END
  END output_thermometer_o[138]
  PIN output_thermometer_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.050 0.000 138.190 0.410 ;
    END
  END output_thermometer_o[48]
  PIN output_binary_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.430 208.350 139.570 210.000 ;
    END
  END output_binary_o[1]
  PIN output_thermometer_o[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.430 0.000 139.570 0.410 ;
    END
  END output_thermometer_o[225]
  PIN output_thermometer_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.810 208.350 140.950 210.000 ;
    END
  END output_thermometer_o[121]
  PIN output_thermometer_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.810 0.000 140.950 0.410 ;
    END
  END output_thermometer_o[10]
  PIN output_thermometer_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.190 208.350 142.330 210.000 ;
    END
  END output_thermometer_o[77]
  PIN output_thermometer_o[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.190 0.000 142.330 1.090 ;
    END
  END output_thermometer_o[170]
  PIN output_thermometer_o[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.570 208.350 143.710 210.000 ;
    END
  END output_thermometer_o[141]
  PIN output_thermometer_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.570 0.000 143.710 0.410 ;
    END
  END output_thermometer_o[40]
  PIN output_thermometer_o[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.950 208.350 145.090 210.000 ;
    END
  END output_thermometer_o[216]
  PIN output_thermometer_o[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.950 0.000 145.090 1.260 ;
    END
  END output_thermometer_o[139]
  PIN output_thermometer_o[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.330 208.350 146.470 210.000 ;
    END
  END output_thermometer_o[210]
  PIN output_thermometer_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.330 0.000 146.470 0.410 ;
    END
  END output_thermometer_o[42]
  PIN output_thermometer_o[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.710 208.350 147.850 210.000 ;
    END
  END output_thermometer_o[150]
  PIN output_thermometer_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.710 0.000 147.850 1.060 ;
    END
  END output_thermometer_o[88]
  PIN output_thermometer_o[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.090 208.350 149.230 210.000 ;
    END
  END output_thermometer_o[240]
  PIN output_thermometer_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.090 0.000 149.230 0.410 ;
    END
  END output_thermometer_o[1]
  PIN output_thermometer_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.470 208.350 150.610 210.000 ;
    END
  END output_thermometer_o[66]
  PIN output_thermometer_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.470 0.000 150.610 0.410 ;
    END
  END output_thermometer_o[36]
  PIN output_thermometer_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.850 208.350 151.990 210.000 ;
    END
  END output_thermometer_o[127]
  PIN output_thermometer_o[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.850 0.000 151.990 0.410 ;
    END
  END output_thermometer_o[177]
  PIN output_thermometer_o[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.230 208.350 153.370 210.000 ;
    END
  END output_thermometer_o[148]
  PIN output_thermometer_o[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.230 0.000 153.370 0.410 ;
    END
  END output_thermometer_o[239]
  PIN output_thermometer_o[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.610 208.350 154.750 210.000 ;
    END
  END output_thermometer_o[255]
  PIN output_thermometer_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.610 0.000 154.750 1.090 ;
    END
  END output_thermometer_o[71]
  PIN output_thermometer_o[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.990 208.350 156.130 210.000 ;
    END
  END output_thermometer_o[133]
  PIN output_thermometer_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.990 0.000 156.130 1.090 ;
    END
  END output_thermometer_o[91]
  PIN output_thermometer_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.370 208.350 157.510 210.000 ;
    END
  END output_thermometer_o[22]
  PIN output_thermometer_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.370 0.000 157.510 1.260 ;
    END
  END output_thermometer_o[65]
  PIN output_thermometer_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.750 208.350 158.890 210.000 ;
    END
  END output_thermometer_o[75]
  PIN output_thermometer_o[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.750 0.000 158.890 0.410 ;
    END
  END output_thermometer_o[192]
  PIN output_thermometer_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.130 208.350 160.270 210.000 ;
    END
  END output_thermometer_o[51]
  PIN output_thermometer_o[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.130 0.000 160.270 0.410 ;
    END
  END output_thermometer_o[171]
  PIN output_thermometer_o[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.510 208.350 161.650 210.000 ;
    END
  END output_thermometer_o[254]
  PIN output_thermometer_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.510 0.000 161.650 0.410 ;
    END
  END output_thermometer_o[28]
  PIN output_thermometer_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.890 208.350 163.030 210.000 ;
    END
  END output_thermometer_o[122]
  PIN output_thermometer_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.890 0.000 163.030 0.410 ;
    END
  END output_thermometer_o[70]
  PIN output_thermometer_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.270 208.350 164.410 210.000 ;
    END
  END output_thermometer_o[46]
  PIN output_thermometer_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.270 0.000 164.410 1.090 ;
    END
  END output_thermometer_o[100]
  PIN output_thermometer_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.650 208.350 165.790 210.000 ;
    END
  END output_thermometer_o[56]
  PIN output_thermometer_o[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.650 0.000 165.790 0.410 ;
    END
  END output_thermometer_o[172]
  PIN output_thermometer_o[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.030 208.350 167.170 210.000 ;
    END
  END output_thermometer_o[135]
  PIN output_thermometer_o[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.030 0.000 167.170 1.260 ;
    END
  END output_thermometer_o[184]
  PIN output_thermometer_o[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.410 208.350 168.550 210.000 ;
    END
  END output_thermometer_o[173]
  PIN output_thermometer_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.410 0.000 168.550 1.090 ;
    END
  END output_thermometer_o[85]
  PIN output_thermometer_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.790 208.350 169.930 210.000 ;
    END
  END output_thermometer_o[38]
  PIN output_thermometer_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.790 0.000 169.930 0.410 ;
    END
  END output_thermometer_o[52]
  PIN output_thermometer_o[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.170 208.350 171.310 210.000 ;
    END
  END output_thermometer_o[238]
  PIN output_thermometer_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.170 0.000 171.310 1.260 ;
    END
  END output_thermometer_o[92]
  PIN output_thermometer_o[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.550 208.350 172.690 210.000 ;
    END
  END output_thermometer_o[165]
  PIN output_thermometer_o[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.550 0.000 172.690 0.410 ;
    END
  END output_thermometer_o[223]
  PIN output_thermometer_o[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.930 208.350 174.070 210.000 ;
    END
  END output_thermometer_o[246]
  PIN output_thermometer_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.930 0.000 174.070 1.090 ;
    END
  END output_thermometer_o[118]
  PIN output_thermometer_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.310 208.350 175.450 210.000 ;
    END
  END output_thermometer_o[50]
  PIN output_thermometer_o[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.310 0.000 175.450 0.410 ;
    END
  END output_thermometer_o[202]
  PIN output_thermometer_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.690 209.030 176.830 210.000 ;
    END
  END output_thermometer_o[113]
  PIN output_thermometer_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.690 0.000 176.830 0.410 ;
    END
  END output_thermometer_o[80]
  PIN output_thermometer_o[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.070 208.350 178.210 210.000 ;
    END
  END output_thermometer_o[231]
  PIN output_thermometer_o[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.070 0.000 178.210 1.260 ;
    END
  END output_thermometer_o[153]
  PIN output_thermometer_o[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.450 208.350 179.590 210.000 ;
    END
  END output_thermometer_o[203]
  PIN output_thermometer_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.450 0.000 179.590 0.410 ;
    END
  END output_thermometer_o[6]
  PIN output_thermometer_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.830 208.350 180.970 210.000 ;
    END
  END output_thermometer_o[44]
  PIN output_thermometer_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.830 0.000 180.970 0.410 ;
    END
  END output_thermometer_o[0]
  PIN output_thermometer_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.210 208.350 182.350 210.000 ;
    END
  END output_thermometer_o[108]
  PIN output_thermometer_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.210 0.000 182.350 0.410 ;
    END
  END output_thermometer_o[24]
  PIN en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.590 208.350 183.730 210.000 ;
    END
  END en_o
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 95.180 270.000 95.780 ;
    END
  END clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 96.540 270.000 97.140 ;
    END
  END rst_ni
  PIN randomise_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 97.900 270.000 98.500 ;
    END
  END randomise_en_i
  PIN en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 99.260 270.000 99.860 ;
    END
  END en_i
  PIN input_binary_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 100.620 270.000 101.220 ;
    END
  END input_binary_i[0]
  PIN input_binary_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 101.980 270.000 102.580 ;
    END
  END input_binary_i[1]
  PIN input_binary_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 103.340 270.000 103.940 ;
    END
  END input_binary_i[2]
  PIN input_binary_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 104.700 270.000 105.300 ;
    END
  END input_binary_i[3]
  PIN input_binary_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 106.060 270.000 106.660 ;
    END
  END input_binary_i[4]
  PIN input_binary_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 107.420 270.000 108.020 ;
    END
  END input_binary_i[5]
  PIN input_binary_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 108.780 270.000 109.380 ;
    END
  END input_binary_i[6]
  PIN input_binary_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 110.140 270.000 110.740 ;
    END
  END input_binary_i[7]
  PIN input_binary_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 111.500 270.000 112.100 ;
    END
  END input_binary_i[8]
  PIN input_binary_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.800 112.860 270.000 113.460 ;
    END
  END input_binary_i[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 198.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 198.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 264.040 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 264.040 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 198.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 198.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 264.040 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 7.905 264.040 205.275 ;
      LAYER met1 ;
        RECT 1.910 0.380 266.270 209.060 ;
      LAYER met2 ;
        RECT 1.940 208.070 5.290 209.170 ;
        RECT 5.990 208.070 6.670 209.170 ;
        RECT 7.370 208.070 8.050 209.170 ;
        RECT 8.750 208.070 9.430 209.170 ;
        RECT 10.130 208.070 10.810 209.170 ;
        RECT 11.510 208.070 12.190 209.170 ;
        RECT 12.890 208.070 13.570 209.170 ;
        RECT 14.270 208.070 14.950 209.170 ;
        RECT 15.650 208.070 16.330 209.170 ;
        RECT 17.030 208.070 17.710 209.170 ;
        RECT 18.410 208.070 19.090 209.170 ;
        RECT 19.790 208.440 20.470 209.170 ;
        RECT 21.170 208.780 21.850 209.170 ;
        RECT 22.550 208.780 23.230 209.170 ;
        RECT 21.170 208.440 23.230 208.780 ;
        RECT 19.790 208.070 23.230 208.440 ;
        RECT 23.930 208.070 24.610 209.170 ;
        RECT 25.310 208.070 25.990 209.170 ;
        RECT 26.690 208.070 27.370 209.170 ;
        RECT 28.070 208.070 28.750 209.170 ;
        RECT 29.450 208.070 30.130 209.170 ;
        RECT 30.830 208.070 31.510 209.170 ;
        RECT 32.210 208.070 32.890 209.170 ;
        RECT 33.590 208.070 34.270 209.170 ;
        RECT 34.970 208.070 35.650 209.170 ;
        RECT 36.350 208.070 37.030 209.170 ;
        RECT 37.730 208.070 38.410 209.170 ;
        RECT 39.110 208.070 39.790 209.170 ;
        RECT 40.490 208.070 41.170 209.170 ;
        RECT 41.870 208.070 42.550 209.170 ;
        RECT 43.250 208.070 43.930 209.170 ;
        RECT 44.630 208.070 45.310 209.170 ;
        RECT 46.010 208.070 46.690 209.170 ;
        RECT 47.390 208.070 48.070 209.170 ;
        RECT 48.770 208.070 49.450 209.170 ;
        RECT 50.150 208.070 50.830 209.170 ;
        RECT 51.530 208.750 52.210 209.170 ;
        RECT 52.910 208.750 53.590 209.170 ;
        RECT 51.530 208.070 53.590 208.750 ;
        RECT 54.290 208.070 54.970 209.170 ;
        RECT 55.670 208.070 56.350 209.170 ;
        RECT 57.050 208.070 57.730 209.170 ;
        RECT 58.430 208.070 59.110 209.170 ;
        RECT 59.810 208.070 60.490 209.170 ;
        RECT 61.190 208.070 61.870 209.170 ;
        RECT 62.570 208.070 63.250 209.170 ;
        RECT 63.950 208.070 64.630 209.170 ;
        RECT 65.330 208.070 66.010 209.170 ;
        RECT 66.710 208.070 67.390 209.170 ;
        RECT 68.090 208.070 68.770 209.170 ;
        RECT 69.470 208.070 70.150 209.170 ;
        RECT 70.850 208.070 71.530 209.170 ;
        RECT 72.230 208.070 72.910 209.170 ;
        RECT 73.610 208.070 74.290 209.170 ;
        RECT 74.990 208.070 75.670 209.170 ;
        RECT 76.370 208.070 77.050 209.170 ;
        RECT 77.750 208.070 78.430 209.170 ;
        RECT 79.130 208.070 79.810 209.170 ;
        RECT 80.510 208.070 81.190 209.170 ;
        RECT 81.890 208.070 82.570 209.170 ;
        RECT 83.270 208.070 83.950 209.170 ;
        RECT 84.650 208.070 85.330 209.170 ;
        RECT 86.030 208.750 86.710 209.170 ;
        RECT 87.410 208.750 88.090 209.170 ;
        RECT 86.030 208.070 88.090 208.750 ;
        RECT 88.790 208.070 89.470 209.170 ;
        RECT 90.170 208.070 90.850 209.170 ;
        RECT 91.550 208.070 92.230 209.170 ;
        RECT 92.930 208.070 93.610 209.170 ;
        RECT 94.310 208.070 94.990 209.170 ;
        RECT 95.690 208.780 96.370 209.170 ;
        RECT 97.070 208.780 97.750 209.170 ;
        RECT 95.690 208.440 97.750 208.780 ;
        RECT 98.450 208.440 99.130 209.170 ;
        RECT 95.690 208.070 99.130 208.440 ;
        RECT 99.830 208.070 100.510 209.170 ;
        RECT 101.210 208.070 101.890 209.170 ;
        RECT 102.590 208.070 103.270 209.170 ;
        RECT 103.970 208.070 104.650 209.170 ;
        RECT 105.350 208.070 106.030 209.170 ;
        RECT 106.730 208.070 107.410 209.170 ;
        RECT 108.110 208.070 108.790 209.170 ;
        RECT 109.490 208.440 110.170 209.170 ;
        RECT 110.870 208.440 111.550 209.170 ;
        RECT 109.490 208.070 111.550 208.440 ;
        RECT 112.250 208.070 112.930 209.170 ;
        RECT 113.630 208.070 114.310 209.170 ;
        RECT 115.010 208.070 115.690 209.170 ;
        RECT 116.390 208.070 117.070 209.170 ;
        RECT 117.770 208.070 118.450 209.170 ;
        RECT 119.150 208.070 119.830 209.170 ;
        RECT 120.530 208.070 121.210 209.170 ;
        RECT 121.910 208.070 122.590 209.170 ;
        RECT 123.290 208.070 123.970 209.170 ;
        RECT 124.670 208.070 125.350 209.170 ;
        RECT 126.050 208.070 126.730 209.170 ;
        RECT 127.430 208.070 128.110 209.170 ;
        RECT 128.810 208.070 129.490 209.170 ;
        RECT 130.190 208.070 130.870 209.170 ;
        RECT 131.570 208.440 132.250 209.170 ;
        RECT 132.950 208.440 133.630 209.170 ;
        RECT 131.570 208.070 133.630 208.440 ;
        RECT 134.330 208.070 135.010 209.170 ;
        RECT 135.710 208.070 136.390 209.170 ;
        RECT 137.090 208.070 137.770 209.170 ;
        RECT 138.470 208.070 139.150 209.170 ;
        RECT 139.850 208.070 140.530 209.170 ;
        RECT 141.230 208.070 141.910 209.170 ;
        RECT 142.610 208.070 143.290 209.170 ;
        RECT 143.990 208.070 144.670 209.170 ;
        RECT 145.370 208.070 146.050 209.170 ;
        RECT 146.750 208.070 147.430 209.170 ;
        RECT 148.130 208.070 148.810 209.170 ;
        RECT 149.510 208.070 150.190 209.170 ;
        RECT 150.890 208.070 151.570 209.170 ;
        RECT 152.270 208.070 152.950 209.170 ;
        RECT 153.650 208.070 154.330 209.170 ;
        RECT 155.030 208.070 155.710 209.170 ;
        RECT 156.410 208.070 157.090 209.170 ;
        RECT 157.790 208.070 158.470 209.170 ;
        RECT 159.170 208.070 159.850 209.170 ;
        RECT 160.550 208.070 161.230 209.170 ;
        RECT 161.930 208.070 162.610 209.170 ;
        RECT 163.310 208.070 163.990 209.170 ;
        RECT 164.690 208.070 165.370 209.170 ;
        RECT 166.070 208.070 166.750 209.170 ;
        RECT 167.450 208.070 168.130 209.170 ;
        RECT 168.830 208.070 169.510 209.170 ;
        RECT 170.210 208.070 170.890 209.170 ;
        RECT 171.590 208.070 172.270 209.170 ;
        RECT 172.970 208.070 173.650 209.170 ;
        RECT 174.350 208.070 175.030 209.170 ;
        RECT 175.730 208.750 176.410 209.170 ;
        RECT 177.110 208.750 177.790 209.170 ;
        RECT 175.730 208.070 177.790 208.750 ;
        RECT 178.490 208.070 179.170 209.170 ;
        RECT 179.870 208.070 180.550 209.170 ;
        RECT 181.250 208.070 181.930 209.170 ;
        RECT 182.630 208.070 183.310 209.170 ;
        RECT 184.010 208.070 266.240 209.170 ;
        RECT 1.940 1.540 266.240 208.070 ;
        RECT 1.940 1.370 78.430 1.540 ;
        RECT 1.940 0.070 5.290 1.370 ;
        RECT 5.990 0.070 6.670 1.370 ;
        RECT 7.370 0.070 8.050 1.370 ;
        RECT 8.750 0.070 9.430 1.370 ;
        RECT 10.130 0.070 10.810 1.370 ;
        RECT 11.510 0.690 13.570 1.370 ;
        RECT 11.510 0.070 12.190 0.690 ;
        RECT 12.890 0.070 13.570 0.690 ;
        RECT 14.270 0.070 14.950 1.370 ;
        RECT 15.650 0.070 16.330 1.370 ;
        RECT 17.030 0.070 17.710 1.370 ;
        RECT 18.410 0.690 25.990 1.370 ;
        RECT 18.410 0.070 19.090 0.690 ;
        RECT 19.790 0.070 20.470 0.690 ;
        RECT 21.170 0.070 21.850 0.690 ;
        RECT 22.550 0.070 23.230 0.690 ;
        RECT 23.930 0.070 24.610 0.690 ;
        RECT 25.310 0.070 25.990 0.690 ;
        RECT 26.690 1.340 28.750 1.370 ;
        RECT 26.690 0.070 27.370 1.340 ;
        RECT 28.070 0.070 28.750 1.340 ;
        RECT 29.450 1.340 32.890 1.370 ;
        RECT 29.450 0.690 31.510 1.340 ;
        RECT 29.450 0.070 30.130 0.690 ;
        RECT 30.830 0.070 31.510 0.690 ;
        RECT 32.210 0.070 32.890 1.340 ;
        RECT 33.590 0.690 38.410 1.370 ;
        RECT 33.590 0.070 34.270 0.690 ;
        RECT 34.970 0.070 35.650 0.690 ;
        RECT 36.350 0.070 37.030 0.690 ;
        RECT 37.730 0.070 38.410 0.690 ;
        RECT 39.110 0.070 39.790 1.370 ;
        RECT 40.490 0.690 46.690 1.370 ;
        RECT 40.490 0.070 41.170 0.690 ;
        RECT 41.870 0.070 42.550 0.690 ;
        RECT 43.250 0.070 43.930 0.690 ;
        RECT 44.630 0.070 45.310 0.690 ;
        RECT 46.010 0.070 46.690 0.690 ;
        RECT 47.390 0.690 54.970 1.370 ;
        RECT 47.390 0.070 48.070 0.690 ;
        RECT 48.770 0.070 49.450 0.690 ;
        RECT 50.150 0.070 50.830 0.690 ;
        RECT 51.530 0.070 52.210 0.690 ;
        RECT 52.910 0.070 53.590 0.690 ;
        RECT 54.290 0.070 54.970 0.690 ;
        RECT 55.670 0.690 59.110 1.370 ;
        RECT 55.670 0.070 56.350 0.690 ;
        RECT 57.050 0.070 57.730 0.690 ;
        RECT 58.430 0.070 59.110 0.690 ;
        RECT 59.810 1.340 66.010 1.370 ;
        RECT 59.810 1.000 63.250 1.340 ;
        RECT 59.810 0.690 61.870 1.000 ;
        RECT 59.810 0.070 60.490 0.690 ;
        RECT 61.190 0.070 61.870 0.690 ;
        RECT 62.570 0.070 63.250 1.000 ;
        RECT 63.950 0.690 66.010 1.340 ;
        RECT 63.950 0.070 64.630 0.690 ;
        RECT 65.330 0.070 66.010 0.690 ;
        RECT 66.710 0.070 67.390 1.370 ;
        RECT 68.090 0.070 68.770 1.370 ;
        RECT 69.470 0.070 70.150 1.370 ;
        RECT 70.850 0.070 71.530 1.370 ;
        RECT 72.230 0.690 78.430 1.370 ;
        RECT 72.230 0.070 72.910 0.690 ;
        RECT 73.610 0.070 74.290 0.690 ;
        RECT 74.990 0.070 75.670 0.690 ;
        RECT 76.370 0.070 77.050 0.690 ;
        RECT 77.750 0.070 78.430 0.690 ;
        RECT 79.130 1.370 97.750 1.540 ;
        RECT 79.130 0.070 79.810 1.370 ;
        RECT 80.510 0.070 81.190 1.370 ;
        RECT 81.890 0.690 85.330 1.370 ;
        RECT 81.890 0.070 82.570 0.690 ;
        RECT 83.270 0.070 83.950 0.690 ;
        RECT 84.650 0.070 85.330 0.690 ;
        RECT 86.030 0.070 86.710 1.370 ;
        RECT 87.410 0.070 88.090 1.370 ;
        RECT 88.790 0.070 89.470 1.370 ;
        RECT 90.170 0.070 90.850 1.370 ;
        RECT 91.550 0.690 94.990 1.370 ;
        RECT 91.550 0.070 92.230 0.690 ;
        RECT 92.930 0.070 93.610 0.690 ;
        RECT 94.310 0.070 94.990 0.690 ;
        RECT 95.690 0.690 97.750 1.370 ;
        RECT 95.690 0.070 96.370 0.690 ;
        RECT 97.070 0.070 97.750 0.690 ;
        RECT 98.450 1.370 106.030 1.540 ;
        RECT 98.450 0.690 104.650 1.370 ;
        RECT 98.450 0.070 99.130 0.690 ;
        RECT 99.830 0.070 100.510 0.690 ;
        RECT 101.210 0.070 101.890 0.690 ;
        RECT 102.590 0.070 103.270 0.690 ;
        RECT 103.970 0.070 104.650 0.690 ;
        RECT 105.350 0.070 106.030 1.370 ;
        RECT 106.730 1.370 114.310 1.540 ;
        RECT 106.730 0.070 107.410 1.370 ;
        RECT 108.110 0.690 111.550 1.370 ;
        RECT 108.110 0.070 108.790 0.690 ;
        RECT 109.490 0.070 110.170 0.690 ;
        RECT 110.870 0.070 111.550 0.690 ;
        RECT 112.250 0.070 112.930 1.370 ;
        RECT 113.630 0.070 114.310 1.370 ;
        RECT 115.010 1.370 144.670 1.540 ;
        RECT 115.010 1.340 121.210 1.370 ;
        RECT 115.010 0.070 115.690 1.340 ;
        RECT 116.390 0.690 121.210 1.340 ;
        RECT 116.390 0.070 117.070 0.690 ;
        RECT 117.770 0.070 118.450 0.690 ;
        RECT 119.150 0.070 119.830 0.690 ;
        RECT 120.530 0.070 121.210 0.690 ;
        RECT 121.910 0.690 123.970 1.370 ;
        RECT 121.910 0.070 122.590 0.690 ;
        RECT 123.290 0.070 123.970 0.690 ;
        RECT 124.670 0.070 125.350 1.370 ;
        RECT 126.050 1.000 129.490 1.370 ;
        RECT 126.050 0.690 128.110 1.000 ;
        RECT 126.050 0.070 126.730 0.690 ;
        RECT 127.430 0.070 128.110 0.690 ;
        RECT 128.810 0.070 129.490 1.000 ;
        RECT 130.190 0.690 132.250 1.370 ;
        RECT 130.190 0.070 130.870 0.690 ;
        RECT 131.570 0.070 132.250 0.690 ;
        RECT 132.950 0.070 133.630 1.370 ;
        RECT 134.330 0.690 141.910 1.370 ;
        RECT 134.330 0.070 135.010 0.690 ;
        RECT 135.710 0.070 136.390 0.690 ;
        RECT 137.090 0.070 137.770 0.690 ;
        RECT 138.470 0.070 139.150 0.690 ;
        RECT 139.850 0.070 140.530 0.690 ;
        RECT 141.230 0.070 141.910 0.690 ;
        RECT 142.610 0.690 144.670 1.370 ;
        RECT 142.610 0.070 143.290 0.690 ;
        RECT 143.990 0.070 144.670 0.690 ;
        RECT 145.370 1.370 157.090 1.540 ;
        RECT 145.370 1.340 154.330 1.370 ;
        RECT 145.370 0.690 147.430 1.340 ;
        RECT 145.370 0.070 146.050 0.690 ;
        RECT 146.750 0.070 147.430 0.690 ;
        RECT 148.130 0.690 154.330 1.340 ;
        RECT 148.130 0.070 148.810 0.690 ;
        RECT 149.510 0.070 150.190 0.690 ;
        RECT 150.890 0.070 151.570 0.690 ;
        RECT 152.270 0.070 152.950 0.690 ;
        RECT 153.650 0.070 154.330 0.690 ;
        RECT 155.030 0.070 155.710 1.370 ;
        RECT 156.410 0.070 157.090 1.370 ;
        RECT 157.790 1.370 166.750 1.540 ;
        RECT 157.790 0.690 163.990 1.370 ;
        RECT 157.790 0.070 158.470 0.690 ;
        RECT 159.170 0.070 159.850 0.690 ;
        RECT 160.550 0.070 161.230 0.690 ;
        RECT 161.930 0.070 162.610 0.690 ;
        RECT 163.310 0.070 163.990 0.690 ;
        RECT 164.690 0.690 166.750 1.370 ;
        RECT 164.690 0.070 165.370 0.690 ;
        RECT 166.070 0.070 166.750 0.690 ;
        RECT 167.450 1.370 170.890 1.540 ;
        RECT 167.450 0.070 168.130 1.370 ;
        RECT 168.830 0.690 170.890 1.370 ;
        RECT 168.830 0.070 169.510 0.690 ;
        RECT 170.210 0.070 170.890 0.690 ;
        RECT 171.590 1.370 177.790 1.540 ;
        RECT 171.590 0.690 173.650 1.370 ;
        RECT 171.590 0.070 172.270 0.690 ;
        RECT 172.970 0.070 173.650 0.690 ;
        RECT 174.350 0.690 177.790 1.370 ;
        RECT 174.350 0.070 175.030 0.690 ;
        RECT 175.730 0.070 176.410 0.690 ;
        RECT 177.110 0.070 177.790 0.690 ;
        RECT 178.490 0.690 266.240 1.540 ;
        RECT 178.490 0.070 179.170 0.690 ;
        RECT 179.870 0.070 180.550 0.690 ;
        RECT 181.250 0.070 181.930 0.690 ;
        RECT 182.630 0.070 266.240 0.690 ;
      LAYER met3 ;
        RECT 2.110 113.860 268.800 206.545 ;
        RECT 2.110 94.780 268.400 113.860 ;
        RECT 2.110 0.175 268.800 94.780 ;
      LAYER met4 ;
        RECT 2.135 199.200 267.425 206.545 ;
        RECT 2.135 10.240 20.640 199.200 ;
        RECT 23.040 10.240 97.440 199.200 ;
        RECT 99.840 10.240 174.240 199.200 ;
        RECT 176.640 10.240 251.040 199.200 ;
        RECT 253.440 10.240 267.425 199.200 ;
        RECT 2.135 0.175 267.425 10.240 ;
      LAYER met5 ;
        RECT 6.100 29.690 242.300 39.900 ;
        RECT 6.100 4.300 242.300 24.890 ;
  END
END dac_digital_interface
END LIBRARY

