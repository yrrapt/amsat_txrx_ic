magic
tech sky130A
magscale 1 2
timestamp 1621163452
<< nwell >>
rect 1066 38885 78882 39451
rect 1066 37797 78882 38363
rect 1066 36709 78882 37275
rect 1066 35621 78882 36187
rect 1066 34533 78882 35099
rect 1066 33445 78882 34011
rect 1066 32357 78882 32923
rect 1066 31269 78882 31835
rect 1066 30181 78882 30747
rect 1066 29093 78882 29659
rect 1066 28005 78882 28571
rect 1066 26917 78882 27483
rect 1066 25829 78882 26395
rect 1066 24741 78882 25307
rect 1066 23653 78882 24219
rect 1066 22565 78882 23131
rect 1066 21477 78882 22043
rect 1066 20389 78882 20955
rect 1066 19301 78882 19867
rect 1066 18213 78882 18779
rect 1066 17125 78882 17691
rect 1066 16037 78882 16603
rect 1066 14949 78882 15515
rect 1066 13861 78882 14427
rect 1066 12773 78882 13339
rect 1066 11685 78882 12251
rect 1066 10597 78882 11163
rect 1066 9509 78882 10075
rect 1066 8421 78882 8987
rect 1066 7333 78882 7899
rect 1066 6245 78882 6811
rect 1066 5157 78882 5723
rect 1066 4069 78882 4635
rect 1066 2981 78882 3547
rect 1066 2138 78882 2459
<< obsli1 >>
rect 1104 1445 78844 41395
<< obsm1 >>
rect 1104 144 79290 41880
<< metal2 >>
rect 1114 41670 1142 42000
rect 1390 41670 1418 42000
rect 1666 41670 1694 42000
rect 1942 41670 1970 42000
rect 2218 41670 2246 42000
rect 2494 41670 2522 42000
rect 2770 41670 2798 42000
rect 3046 41670 3074 42000
rect 3322 41670 3350 42000
rect 3598 41670 3626 42000
rect 3874 41670 3902 42000
rect 4150 41670 4178 42000
rect 4426 41670 4454 42000
rect 4702 41806 4730 42000
rect 4978 41670 5006 42000
rect 5254 41670 5282 42000
rect 5530 41670 5558 42000
rect 5806 41670 5834 42000
rect 6082 41670 6110 42000
rect 6358 41744 6386 42000
rect 6634 41670 6662 42000
rect 6910 41670 6938 42000
rect 7186 41670 7214 42000
rect 7462 41670 7490 42000
rect 7738 41670 7766 42000
rect 8014 41670 8042 42000
rect 8290 41670 8318 42000
rect 8566 41670 8594 42000
rect 8842 41670 8870 42000
rect 9118 41670 9146 42000
rect 9394 41670 9422 42000
rect 9670 41670 9698 42000
rect 9946 41670 9974 42000
rect 10222 41670 10250 42000
rect 10498 41670 10526 42000
rect 10774 41670 10802 42000
rect 11050 41744 11078 42000
rect 11326 41670 11354 42000
rect 11602 41670 11630 42000
rect 11878 41670 11906 42000
rect 12154 41670 12182 42000
rect 12430 41670 12458 42000
rect 12706 41670 12734 42000
rect 12982 41670 13010 42000
rect 13258 41670 13286 42000
rect 13534 41670 13562 42000
rect 13810 41670 13838 42000
rect 14086 41670 14114 42000
rect 14362 41670 14390 42000
rect 14638 41670 14666 42000
rect 14914 41670 14942 42000
rect 15190 41670 15218 42000
rect 15466 41806 15494 42000
rect 15742 41670 15770 42000
rect 16018 41670 16046 42000
rect 16294 41744 16322 42000
rect 16570 41670 16598 42000
rect 16846 41670 16874 42000
rect 17122 41670 17150 42000
rect 17398 41670 17426 42000
rect 17674 41670 17702 42000
rect 17950 41670 17978 42000
rect 18226 41670 18254 42000
rect 18502 41670 18530 42000
rect 18778 41670 18806 42000
rect 19054 41670 19082 42000
rect 19330 41744 19358 42000
rect 19606 41670 19634 42000
rect 19882 41670 19910 42000
rect 20158 41670 20186 42000
rect 20434 41670 20462 42000
rect 20710 41670 20738 42000
rect 20986 41670 21014 42000
rect 21262 41806 21290 42000
rect 21538 41670 21566 42000
rect 21814 41806 21842 42000
rect 22090 41670 22118 42000
rect 22366 41670 22394 42000
rect 22642 41670 22670 42000
rect 22918 41670 22946 42000
rect 23194 41670 23222 42000
rect 23470 41670 23498 42000
rect 23746 41670 23774 42000
rect 24022 41670 24050 42000
rect 24298 41670 24326 42000
rect 24574 41670 24602 42000
rect 24850 41670 24878 42000
rect 25126 41670 25154 42000
rect 25402 41670 25430 42000
rect 25678 41670 25706 42000
rect 25954 41670 25982 42000
rect 26230 41670 26258 42000
rect 26506 41670 26534 42000
rect 26782 41670 26810 42000
rect 27058 41670 27086 42000
rect 27334 41670 27362 42000
rect 27610 41670 27638 42000
rect 27886 41670 27914 42000
rect 28162 41670 28190 42000
rect 28438 41670 28466 42000
rect 28714 41670 28742 42000
rect 28990 41670 29018 42000
rect 29266 41670 29294 42000
rect 29542 41670 29570 42000
rect 29818 41744 29846 42000
rect 30094 41670 30122 42000
rect 30370 41670 30398 42000
rect 30646 41670 30674 42000
rect 30922 41670 30950 42000
rect 31198 41670 31226 42000
rect 31474 41670 31502 42000
rect 31750 41880 31778 42000
rect 32026 41670 32054 42000
rect 32302 41670 32330 42000
rect 32578 41670 32606 42000
rect 32854 41670 32882 42000
rect 33130 41744 33158 42000
rect 33406 41806 33434 42000
rect 33682 41812 33710 42000
rect 33958 41670 33986 42000
rect 34234 41670 34262 42000
rect 34510 41670 34538 42000
rect 34786 41670 34814 42000
rect 35062 41670 35090 42000
rect 35338 41806 35366 42000
rect 35614 41670 35642 42000
rect 35890 41670 35918 42000
rect 36166 41670 36194 42000
rect 36442 41744 36470 42000
rect 36718 41670 36746 42000
rect 1114 0 1142 218
rect 1390 0 1418 82
rect 1666 0 1694 218
rect 1942 0 1970 82
rect 2218 0 2246 218
rect 2494 0 2522 218
rect 2770 0 2798 82
rect 3046 0 3074 82
rect 3322 0 3350 218
rect 3598 0 3626 218
rect 3874 0 3902 218
rect 4150 0 4178 82
rect 4426 0 4454 82
rect 4702 0 4730 218
rect 4978 0 5006 82
rect 5254 0 5282 82
rect 5530 0 5558 82
rect 5806 0 5834 82
rect 6082 0 6110 218
rect 6358 0 6386 82
rect 6634 0 6662 82
rect 6910 0 6938 82
rect 7186 0 7214 82
rect 7462 0 7490 218
rect 7738 0 7766 218
rect 8014 0 8042 218
rect 8290 0 8318 218
rect 8566 0 8594 82
rect 8842 0 8870 82
rect 9118 0 9146 82
rect 9394 0 9422 218
rect 9670 0 9698 218
rect 9946 0 9974 218
rect 10222 0 10250 212
rect 10498 0 10526 218
rect 10774 0 10802 82
rect 11050 0 11078 82
rect 11326 0 11354 82
rect 11602 0 11630 218
rect 11878 0 11906 82
rect 12154 0 12182 218
rect 12430 0 12458 82
rect 12706 0 12734 218
rect 12982 0 13010 218
rect 13258 0 13286 218
rect 13534 0 13562 82
rect 13810 0 13838 218
rect 14086 0 14114 82
rect 14362 0 14390 82
rect 14638 0 14666 82
rect 14914 0 14942 144
rect 15190 0 15218 212
rect 15466 0 15494 218
rect 15742 0 15770 218
rect 16018 0 16046 218
rect 16294 0 16322 82
rect 16570 0 16598 218
rect 16846 0 16874 82
rect 17122 0 17150 82
rect 17398 0 17426 82
rect 17674 0 17702 82
rect 17950 0 17978 218
rect 18226 0 18254 82
rect 18502 0 18530 82
rect 18778 0 18806 218
rect 19054 0 19082 82
rect 19330 0 19358 144
rect 19606 0 19634 82
rect 19882 0 19910 82
rect 20158 0 20186 82
rect 20434 0 20462 82
rect 20710 0 20738 218
rect 20986 0 21014 218
rect 21262 0 21290 82
rect 21538 0 21566 82
rect 21814 0 21842 218
rect 22090 0 22118 218
rect 22366 0 22394 218
rect 22642 0 22670 82
rect 22918 0 22946 82
rect 23194 0 23222 82
rect 23470 0 23498 82
rect 23746 0 23774 218
rect 24022 0 24050 82
rect 24298 0 24326 82
rect 24574 0 24602 218
rect 24850 0 24878 218
rect 25126 0 25154 218
rect 25402 0 25430 218
rect 25678 0 25706 212
rect 25954 0 25982 252
rect 26230 0 26258 82
rect 26506 0 26534 218
rect 26782 0 26810 218
rect 27058 0 27086 82
rect 27334 0 27362 218
rect 27610 0 27638 82
rect 27886 0 27914 82
rect 28162 0 28190 218
rect 28438 0 28466 82
rect 28714 0 28742 82
rect 28990 0 29018 82
rect 29266 0 29294 82
rect 29542 0 29570 252
rect 29818 0 29846 82
rect 30094 0 30122 218
rect 30370 0 30398 82
rect 30646 0 30674 82
rect 30922 0 30950 82
rect 31198 0 31226 82
rect 31474 0 31502 218
rect 31750 0 31778 82
rect 32026 0 32054 218
rect 32302 0 32330 82
rect 32578 0 32606 82
rect 32854 0 32882 218
rect 33130 0 33158 212
rect 33406 0 33434 82
rect 33682 0 33710 82
rect 33958 0 33986 218
rect 34234 0 34262 82
rect 34510 0 34538 82
rect 34786 0 34814 218
rect 35062 0 35090 82
rect 35338 0 35366 218
rect 35614 0 35642 218
rect 35890 0 35918 82
rect 36166 0 36194 218
rect 36442 0 36470 218
<< obsm2 >>
rect 1198 41614 1334 41886
rect 1474 41614 1610 41886
rect 1750 41614 1886 41886
rect 2026 41614 2162 41886
rect 2302 41614 2438 41886
rect 2578 41614 2714 41886
rect 2854 41614 2990 41886
rect 3130 41614 3266 41886
rect 3406 41614 3542 41886
rect 3682 41614 3818 41886
rect 3958 41614 4094 41886
rect 4234 41614 4370 41886
rect 4510 41750 4646 41886
rect 4786 41750 4922 41886
rect 4510 41614 4922 41750
rect 5062 41614 5198 41886
rect 5338 41614 5474 41886
rect 5614 41614 5750 41886
rect 5890 41614 6026 41886
rect 6166 41688 6302 41886
rect 6442 41688 6578 41886
rect 6166 41614 6578 41688
rect 6718 41614 6854 41886
rect 6994 41614 7130 41886
rect 7270 41614 7406 41886
rect 7546 41614 7682 41886
rect 7822 41614 7958 41886
rect 8098 41614 8234 41886
rect 8374 41614 8510 41886
rect 8650 41614 8786 41886
rect 8926 41614 9062 41886
rect 9202 41614 9338 41886
rect 9478 41614 9614 41886
rect 9754 41614 9890 41886
rect 10030 41614 10166 41886
rect 10306 41614 10442 41886
rect 10582 41614 10718 41886
rect 10858 41688 10994 41886
rect 11134 41688 11270 41886
rect 10858 41614 11270 41688
rect 11410 41614 11546 41886
rect 11686 41614 11822 41886
rect 11962 41614 12098 41886
rect 12238 41614 12374 41886
rect 12514 41614 12650 41886
rect 12790 41614 12926 41886
rect 13066 41614 13202 41886
rect 13342 41614 13478 41886
rect 13618 41614 13754 41886
rect 13894 41614 14030 41886
rect 14170 41614 14306 41886
rect 14446 41614 14582 41886
rect 14722 41614 14858 41886
rect 14998 41614 15134 41886
rect 15274 41750 15410 41886
rect 15550 41750 15686 41886
rect 15274 41614 15686 41750
rect 15826 41614 15962 41886
rect 16102 41688 16238 41886
rect 16378 41688 16514 41886
rect 16102 41614 16514 41688
rect 16654 41614 16790 41886
rect 16930 41614 17066 41886
rect 17206 41614 17342 41886
rect 17482 41614 17618 41886
rect 17758 41614 17894 41886
rect 18034 41614 18170 41886
rect 18310 41614 18446 41886
rect 18586 41614 18722 41886
rect 18862 41614 18998 41886
rect 19138 41688 19274 41886
rect 19414 41688 19550 41886
rect 19138 41614 19550 41688
rect 19690 41614 19826 41886
rect 19966 41614 20102 41886
rect 20242 41614 20378 41886
rect 20518 41614 20654 41886
rect 20794 41614 20930 41886
rect 21070 41750 21206 41886
rect 21346 41750 21482 41886
rect 21070 41614 21482 41750
rect 21622 41750 21758 41886
rect 21898 41750 22034 41886
rect 21622 41614 22034 41750
rect 22174 41614 22310 41886
rect 22450 41614 22586 41886
rect 22726 41614 22862 41886
rect 23002 41614 23138 41886
rect 23278 41614 23414 41886
rect 23554 41614 23690 41886
rect 23830 41614 23966 41886
rect 24106 41614 24242 41886
rect 24382 41614 24518 41886
rect 24658 41614 24794 41886
rect 24934 41614 25070 41886
rect 25210 41614 25346 41886
rect 25486 41614 25622 41886
rect 25762 41614 25898 41886
rect 26038 41614 26174 41886
rect 26314 41614 26450 41886
rect 26590 41614 26726 41886
rect 26866 41614 27002 41886
rect 27142 41614 27278 41886
rect 27418 41614 27554 41886
rect 27694 41614 27830 41886
rect 27970 41614 28106 41886
rect 28246 41614 28382 41886
rect 28522 41614 28658 41886
rect 28798 41614 28934 41886
rect 29074 41614 29210 41886
rect 29350 41614 29486 41886
rect 29626 41688 29762 41886
rect 29902 41688 30038 41886
rect 29626 41614 30038 41688
rect 30178 41614 30314 41886
rect 30454 41614 30590 41886
rect 30730 41614 30866 41886
rect 31006 41614 31142 41886
rect 31282 41614 31418 41886
rect 31558 41824 31694 41886
rect 31834 41824 31970 41886
rect 31558 41614 31970 41824
rect 32110 41614 32246 41886
rect 32386 41614 32522 41886
rect 32662 41614 32798 41886
rect 32938 41688 33074 41886
rect 33214 41750 33350 41886
rect 33490 41756 33626 41886
rect 33766 41756 33902 41886
rect 33490 41750 33902 41756
rect 33214 41688 33902 41750
rect 32938 41614 33902 41688
rect 34042 41614 34178 41886
rect 34318 41614 34454 41886
rect 34594 41614 34730 41886
rect 34870 41614 35006 41886
rect 35146 41750 35282 41886
rect 35422 41750 35558 41886
rect 35146 41614 35558 41750
rect 35698 41614 35834 41886
rect 35974 41614 36110 41886
rect 36250 41688 36386 41886
rect 36526 41688 36662 41886
rect 36250 41614 36662 41688
rect 36802 41614 79286 41886
rect 1124 308 79286 41614
rect 1124 274 25898 308
rect 1198 138 1610 274
rect 1198 14 1334 138
rect 1474 14 1610 138
rect 1750 138 2162 274
rect 1750 14 1886 138
rect 2026 14 2162 138
rect 2302 14 2438 274
rect 2578 138 3266 274
rect 2578 14 2714 138
rect 2854 14 2990 138
rect 3130 14 3266 138
rect 3406 14 3542 274
rect 3682 14 3818 274
rect 3958 138 4646 274
rect 3958 14 4094 138
rect 4234 14 4370 138
rect 4510 14 4646 138
rect 4786 138 6026 274
rect 4786 14 4922 138
rect 5062 14 5198 138
rect 5338 14 5474 138
rect 5614 14 5750 138
rect 5890 14 6026 138
rect 6166 138 7406 274
rect 6166 14 6302 138
rect 6442 14 6578 138
rect 6718 14 6854 138
rect 6994 14 7130 138
rect 7270 14 7406 138
rect 7546 14 7682 274
rect 7822 14 7958 274
rect 8098 14 8234 274
rect 8374 138 9338 274
rect 8374 14 8510 138
rect 8650 14 8786 138
rect 8926 14 9062 138
rect 9202 14 9338 138
rect 9478 14 9614 274
rect 9754 14 9890 274
rect 10030 268 10442 274
rect 10030 14 10166 268
rect 10306 14 10442 268
rect 10582 138 11546 274
rect 10582 14 10718 138
rect 10858 14 10994 138
rect 11134 14 11270 138
rect 11410 14 11546 138
rect 11686 138 12098 274
rect 11686 14 11822 138
rect 11962 14 12098 138
rect 12238 138 12650 274
rect 12238 14 12374 138
rect 12514 14 12650 138
rect 12790 14 12926 274
rect 13066 14 13202 274
rect 13342 138 13754 274
rect 13894 268 15410 274
rect 13342 14 13478 138
rect 13618 14 13754 138
rect 13894 200 15134 268
rect 13894 138 14858 200
rect 13894 14 14030 138
rect 14170 14 14306 138
rect 14446 14 14582 138
rect 14722 14 14858 138
rect 14998 14 15134 200
rect 15274 14 15410 268
rect 15550 14 15686 274
rect 15826 14 15962 274
rect 16102 138 16514 274
rect 16102 14 16238 138
rect 16378 14 16514 138
rect 16654 138 17894 274
rect 16654 14 16790 138
rect 16930 14 17066 138
rect 17206 14 17342 138
rect 17482 14 17618 138
rect 17758 14 17894 138
rect 18034 138 18722 274
rect 18034 14 18170 138
rect 18310 14 18446 138
rect 18586 14 18722 138
rect 18862 200 20654 274
rect 18862 138 19274 200
rect 18862 14 18998 138
rect 19138 14 19274 138
rect 19414 138 20654 200
rect 19414 14 19550 138
rect 19690 14 19826 138
rect 19966 14 20102 138
rect 20242 14 20378 138
rect 20518 14 20654 138
rect 20794 14 20930 274
rect 21070 138 21758 274
rect 21070 14 21206 138
rect 21346 14 21482 138
rect 21622 14 21758 138
rect 21898 14 22034 274
rect 22174 14 22310 274
rect 22450 138 23690 274
rect 22450 14 22586 138
rect 22726 14 22862 138
rect 23002 14 23138 138
rect 23278 14 23414 138
rect 23554 14 23690 138
rect 23830 138 24518 274
rect 23830 14 23966 138
rect 24106 14 24242 138
rect 24382 14 24518 138
rect 24658 14 24794 274
rect 24934 14 25070 274
rect 25210 14 25346 274
rect 25486 268 25898 274
rect 25486 14 25622 268
rect 25762 14 25898 268
rect 26038 274 29486 308
rect 26038 138 26450 274
rect 26038 14 26174 138
rect 26314 14 26450 138
rect 26590 14 26726 274
rect 26866 138 27278 274
rect 26866 14 27002 138
rect 27142 14 27278 138
rect 27418 138 28106 274
rect 27418 14 27554 138
rect 27694 14 27830 138
rect 27970 14 28106 138
rect 28246 138 29486 274
rect 29626 274 79286 308
rect 28246 14 28382 138
rect 28522 14 28658 138
rect 28798 14 28934 138
rect 29074 14 29210 138
rect 29350 14 29486 138
rect 29626 138 30038 274
rect 29626 14 29762 138
rect 29902 14 30038 138
rect 30178 138 31418 274
rect 30178 14 30314 138
rect 30454 14 30590 138
rect 30730 14 30866 138
rect 31006 14 31142 138
rect 31282 14 31418 138
rect 31558 138 31970 274
rect 31558 14 31694 138
rect 31834 14 31970 138
rect 32110 138 32798 274
rect 32938 268 33902 274
rect 32110 14 32246 138
rect 32386 14 32522 138
rect 32662 14 32798 138
rect 32938 14 33074 268
rect 33214 138 33902 268
rect 33214 14 33350 138
rect 33490 14 33626 138
rect 33766 14 33902 138
rect 34042 138 34730 274
rect 34042 14 34178 138
rect 34318 14 34454 138
rect 34594 14 34730 138
rect 34870 138 35282 274
rect 34870 14 35006 138
rect 35146 14 35282 138
rect 35422 14 35558 274
rect 35698 138 36110 274
rect 35698 14 35834 138
rect 35974 14 36110 138
rect 36250 14 36386 274
rect 36526 14 79286 274
<< metal3 >>
rect 79760 22572 80000 22692
rect 79760 22300 80000 22420
rect 79760 22028 80000 22148
rect 79760 21756 80000 21876
rect 79760 21484 80000 21604
rect 79760 21212 80000 21332
rect 79760 20940 80000 21060
rect 79760 20668 80000 20788
rect 79760 20396 80000 20516
rect 79760 20124 80000 20244
rect 79760 19852 80000 19972
rect 79760 19580 80000 19700
rect 79760 19308 80000 19428
rect 79760 19036 80000 19156
<< obsm3 >>
rect 2681 22772 79760 40357
rect 2681 18956 79680 22772
rect 2681 171 79760 18956
<< metal4 >>
rect 4208 2128 4528 39760
rect 19568 2128 19888 39760
rect 34928 2128 35248 39760
rect 50288 2128 50608 39760
rect 65648 2128 65968 39760
<< obsm4 >>
rect 8070 2048 19488 36821
rect 19968 2048 34848 36821
rect 35328 2048 50208 36821
rect 50688 2048 65568 36821
rect 66048 2048 66181 36821
rect 8070 902 66181 2048
<< metal5 >>
rect 1104 35934 78844 36254
rect 1104 20616 78844 20936
rect 1104 5298 78844 5618
<< obsm5 >>
rect 8028 860 58028 1180
<< labels >>
rlabel metal2 s 1114 41670 1142 42000 6 output_thermometer_o[69]
port 1 nsew signal output
rlabel metal2 s 1114 0 1142 218 6 output_thermometer_o[112]
port 2 nsew signal output
rlabel metal2 s 1390 41670 1418 42000 6 output_thermometer_o[244]
port 3 nsew signal output
rlabel metal2 s 1390 0 1418 82 6 output_thermometer_o[83]
port 4 nsew signal output
rlabel metal2 s 1666 41670 1694 42000 6 output_thermometer_o[54]
port 5 nsew signal output
rlabel metal2 s 1666 0 1694 218 6 output_thermometer_o[166]
port 6 nsew signal output
rlabel metal2 s 1942 41670 1970 42000 6 output_thermometer_o[200]
port 7 nsew signal output
rlabel metal2 s 1942 0 1970 82 6 output_thermometer_o[17]
port 8 nsew signal output
rlabel metal2 s 2218 41670 2246 42000 6 output_thermometer_o[195]
port 9 nsew signal output
rlabel metal2 s 2218 0 2246 218 6 output_thermometer_o[15]
port 10 nsew signal output
rlabel metal2 s 2494 41670 2522 42000 6 output_thermometer_o[130]
port 11 nsew signal output
rlabel metal2 s 2494 0 2522 218 6 output_thermometer_o[229]
port 12 nsew signal output
rlabel metal2 s 2770 41670 2798 42000 6 output_thermometer_o[82]
port 13 nsew signal output
rlabel metal2 s 2770 0 2798 82 6 output_thermometer_o[4]
port 14 nsew signal output
rlabel metal2 s 3046 41670 3074 42000 6 output_thermometer_o[245]
port 15 nsew signal output
rlabel metal2 s 3046 0 3074 82 6 output_thermometer_o[61]
port 16 nsew signal output
rlabel metal2 s 3322 41670 3350 42000 6 output_thermometer_o[197]
port 17 nsew signal output
rlabel metal2 s 3322 0 3350 218 6 output_thermometer_o[101]
port 18 nsew signal output
rlabel metal2 s 3598 41670 3626 42000 6 output_thermometer_o[251]
port 19 nsew signal output
rlabel metal2 s 3598 0 3626 218 6 output_thermometer_o[213]
port 20 nsew signal output
rlabel metal2 s 3874 41670 3902 42000 6 output_thermometer_o[72]
port 21 nsew signal output
rlabel metal2 s 3874 0 3902 218 6 output_thermometer_o[43]
port 22 nsew signal output
rlabel metal2 s 4150 41670 4178 42000 6 output_thermometer_o[230]
port 23 nsew signal output
rlabel metal2 s 4150 0 4178 82 6 output_thermometer_o[134]
port 24 nsew signal output
rlabel metal2 s 4426 41670 4454 42000 6 output_thermometer_o[115]
port 25 nsew signal output
rlabel metal2 s 4426 0 4454 82 6 output_thermometer_o[212]
port 26 nsew signal output
rlabel metal2 s 4702 41806 4730 42000 6 output_thermometer_o[151]
port 27 nsew signal output
rlabel metal2 s 4702 0 4730 218 6 output_thermometer_o[236]
port 28 nsew signal output
rlabel metal2 s 4978 41670 5006 42000 6 output_thermometer_o[105]
port 29 nsew signal output
rlabel metal2 s 4978 0 5006 82 6 output_thermometer_o[174]
port 30 nsew signal output
rlabel metal2 s 5254 41670 5282 42000 6 output_thermometer_o[196]
port 31 nsew signal output
rlabel metal2 s 5254 0 5282 82 6 output_thermometer_o[57]
port 32 nsew signal output
rlabel metal2 s 5530 41670 5558 42000 6 output_thermometer_o[76]
port 33 nsew signal output
rlabel metal2 s 5530 0 5558 82 6 output_thermometer_o[142]
port 34 nsew signal output
rlabel metal2 s 5806 41670 5834 42000 6 output_thermometer_o[241]
port 35 nsew signal output
rlabel metal2 s 5806 0 5834 82 6 output_thermometer_o[110]
port 36 nsew signal output
rlabel metal2 s 6082 41670 6110 42000 6 output_thermometer_o[123]
port 37 nsew signal output
rlabel metal2 s 6082 0 6110 218 6 output_thermometer_o[81]
port 38 nsew signal output
rlabel metal2 s 6358 41744 6386 42000 6 output_thermometer_o[242]
port 39 nsew signal output
rlabel metal2 s 6358 0 6386 82 6 output_thermometer_o[14]
port 40 nsew signal output
rlabel metal2 s 6634 41670 6662 42000 6 output_thermometer_o[218]
port 41 nsew signal output
rlabel metal2 s 6634 0 6662 82 6 output_thermometer_o[250]
port 42 nsew signal output
rlabel metal2 s 6910 41670 6938 42000 6 output_thermometer_o[94]
port 43 nsew signal output
rlabel metal2 s 6910 0 6938 82 6 output_thermometer_o[129]
port 44 nsew signal output
rlabel metal2 s 7186 41670 7214 42000 6 output_thermometer_o[9]
port 45 nsew signal output
rlabel metal2 s 7186 0 7214 82 6 output_thermometer_o[117]
port 46 nsew signal output
rlabel metal2 s 7462 41670 7490 42000 6 output_thermometer_o[179]
port 47 nsew signal output
rlabel metal2 s 7462 0 7490 218 6 output_thermometer_o[73]
port 48 nsew signal output
rlabel metal2 s 7738 41670 7766 42000 6 output_thermometer_o[86]
port 49 nsew signal output
rlabel metal2 s 7738 0 7766 218 6 output_thermometer_o[215]
port 50 nsew signal output
rlabel metal2 s 8014 41670 8042 42000 6 output_thermometer_o[182]
port 51 nsew signal output
rlabel metal2 s 8014 0 8042 218 6 output_thermometer_o[12]
port 52 nsew signal output
rlabel metal2 s 8290 41670 8318 42000 6 output_thermometer_o[96]
port 53 nsew signal output
rlabel metal2 s 8290 0 8318 218 6 output_thermometer_o[132]
port 54 nsew signal output
rlabel metal2 s 8566 41670 8594 42000 6 output_thermometer_o[29]
port 55 nsew signal output
rlabel metal2 s 8566 0 8594 82 6 output_thermometer_o[232]
port 56 nsew signal output
rlabel metal2 s 8842 41670 8870 42000 6 output_thermometer_o[191]
port 57 nsew signal output
rlabel metal2 s 8842 0 8870 82 6 output_thermometer_o[5]
port 58 nsew signal output
rlabel metal2 s 9118 41670 9146 42000 6 output_thermometer_o[33]
port 59 nsew signal output
rlabel metal2 s 9118 0 9146 82 6 output_thermometer_o[161]
port 60 nsew signal output
rlabel metal2 s 9394 41670 9422 42000 6 output_thermometer_o[11]
port 61 nsew signal output
rlabel metal2 s 9394 0 9422 218 6 output_thermometer_o[160]
port 62 nsew signal output
rlabel metal2 s 9670 41670 9698 42000 6 output_thermometer_o[208]
port 63 nsew signal output
rlabel metal2 s 9670 0 9698 218 6 output_thermometer_o[47]
port 64 nsew signal output
rlabel metal2 s 9946 41670 9974 42000 6 output_thermometer_o[187]
port 65 nsew signal output
rlabel metal2 s 9946 0 9974 218 6 output_thermometer_o[79]
port 66 nsew signal output
rlabel metal2 s 10222 41670 10250 42000 6 output_thermometer_o[59]
port 67 nsew signal output
rlabel metal2 s 10222 0 10250 212 6 output_thermometer_o[116]
port 68 nsew signal output
rlabel metal2 s 10498 41670 10526 42000 6 output_thermometer_o[30]
port 69 nsew signal output
rlabel metal2 s 10498 0 10526 218 6 output_thermometer_o[194]
port 70 nsew signal output
rlabel metal2 s 10774 41670 10802 42000 6 output_thermometer_o[235]
port 71 nsew signal output
rlabel metal2 s 10774 0 10802 82 6 output_thermometer_o[227]
port 72 nsew signal output
rlabel metal2 s 11050 41744 11078 42000 6 output_thermometer_o[97]
port 73 nsew signal output
rlabel metal2 s 11050 0 11078 82 6 output_thermometer_o[67]
port 74 nsew signal output
rlabel metal2 s 11326 41670 11354 42000 6 output_thermometer_o[188]
port 75 nsew signal output
rlabel metal2 s 11326 0 11354 82 6 output_thermometer_o[31]
port 76 nsew signal output
rlabel metal2 s 11602 41670 11630 42000 6 output_thermometer_o[185]
port 77 nsew signal output
rlabel metal2 s 11602 0 11630 218 6 output_thermometer_o[20]
port 78 nsew signal output
rlabel metal2 s 11878 41670 11906 42000 6 output_thermometer_o[32]
port 79 nsew signal output
rlabel metal2 s 11878 0 11906 82 6 output_thermometer_o[125]
port 80 nsew signal output
rlabel metal2 s 12154 41670 12182 42000 6 output_thermometer_o[7]
port 81 nsew signal output
rlabel metal2 s 12154 0 12182 218 6 output_thermometer_o[21]
port 82 nsew signal output
rlabel metal2 s 12430 41670 12458 42000 6 output_thermometer_o[221]
port 83 nsew signal output
rlabel metal2 s 12430 0 12458 82 6 output_thermometer_o[190]
port 84 nsew signal output
rlabel metal2 s 12706 41670 12734 42000 6 output_thermometer_o[37]
port 85 nsew signal output
rlabel metal2 s 12706 0 12734 218 6 output_thermometer_o[74]
port 86 nsew signal output
rlabel metal2 s 12982 41670 13010 42000 6 output_thermometer_o[211]
port 87 nsew signal output
rlabel metal2 s 12982 0 13010 218 6 output_thermometer_o[198]
port 88 nsew signal output
rlabel metal2 s 13258 41670 13286 42000 6 output_thermometer_o[226]
port 89 nsew signal output
rlabel metal2 s 13258 0 13286 218 6 output_thermometer_o[193]
port 90 nsew signal output
rlabel metal2 s 13534 41670 13562 42000 6 output_thermometer_o[249]
port 91 nsew signal output
rlabel metal2 s 13534 0 13562 82 6 output_thermometer_o[84]
port 92 nsew signal output
rlabel metal2 s 13810 41670 13838 42000 6 output_thermometer_o[109]
port 93 nsew signal output
rlabel metal2 s 13810 0 13838 218 6 output_thermometer_o[253]
port 94 nsew signal output
rlabel metal2 s 14086 41670 14114 42000 6 output_thermometer_o[60]
port 95 nsew signal output
rlabel metal2 s 14086 0 14114 82 6 output_thermometer_o[64]
port 96 nsew signal output
rlabel metal2 s 14362 41670 14390 42000 6 output_thermometer_o[23]
port 97 nsew signal output
rlabel metal2 s 14362 0 14390 82 6 output_thermometer_o[164]
port 98 nsew signal output
rlabel metal2 s 14638 41670 14666 42000 6 output_thermometer_o[243]
port 99 nsew signal output
rlabel metal2 s 14638 0 14666 82 6 output_thermometer_o[137]
port 100 nsew signal output
rlabel metal2 s 14914 41670 14942 42000 6 output_thermometer_o[157]
port 101 nsew signal output
rlabel metal2 s 14914 0 14942 144 6 output_thermometer_o[119]
port 102 nsew signal output
rlabel metal2 s 15190 41670 15218 42000 6 output_thermometer_o[217]
port 103 nsew signal output
rlabel metal2 s 15190 0 15218 212 6 output_thermometer_o[90]
port 104 nsew signal output
rlabel metal2 s 15466 41806 15494 42000 6 output_thermometer_o[163]
port 105 nsew signal output
rlabel metal2 s 15466 0 15494 218 6 output_thermometer_o[18]
port 106 nsew signal output
rlabel metal2 s 15742 41670 15770 42000 6 output_thermometer_o[93]
port 107 nsew signal output
rlabel metal2 s 15742 0 15770 218 6 output_thermometer_o[26]
port 108 nsew signal output
rlabel metal2 s 16018 41670 16046 42000 6 output_thermometer_o[107]
port 109 nsew signal output
rlabel metal2 s 16018 0 16046 218 6 output_thermometer_o[144]
port 110 nsew signal output
rlabel metal2 s 16294 41744 16322 42000 6 output_thermometer_o[27]
port 111 nsew signal output
rlabel metal2 s 16294 0 16322 82 6 output_thermometer_o[201]
port 112 nsew signal output
rlabel metal2 s 16570 41670 16598 42000 6 output_thermometer_o[162]
port 113 nsew signal output
rlabel metal2 s 16570 0 16598 218 6 output_thermometer_o[146]
port 114 nsew signal output
rlabel metal2 s 16846 41670 16874 42000 6 output_thermometer_o[168]
port 115 nsew signal output
rlabel metal2 s 16846 0 16874 82 6 output_thermometer_o[53]
port 116 nsew signal output
rlabel metal2 s 17122 41670 17150 42000 6 output_thermometer_o[199]
port 117 nsew signal output
rlabel metal2 s 17122 0 17150 82 6 output_thermometer_o[147]
port 118 nsew signal output
rlabel metal2 s 17398 41670 17426 42000 6 output_thermometer_o[2]
port 119 nsew signal output
rlabel metal2 s 17398 0 17426 82 6 output_thermometer_o[3]
port 120 nsew signal output
rlabel metal2 s 17674 41670 17702 42000 6 output_thermometer_o[136]
port 121 nsew signal output
rlabel metal2 s 17674 0 17702 82 6 output_thermometer_o[204]
port 122 nsew signal output
rlabel metal2 s 17950 41670 17978 42000 6 output_thermometer_o[8]
port 123 nsew signal output
rlabel metal2 s 17950 0 17978 218 6 output_thermometer_o[102]
port 124 nsew signal output
rlabel metal2 s 18226 41670 18254 42000 6 output_thermometer_o[209]
port 125 nsew signal output
rlabel metal2 s 18226 0 18254 82 6 output_thermometer_o[234]
port 126 nsew signal output
rlabel metal2 s 18502 41670 18530 42000 6 output_thermometer_o[145]
port 127 nsew signal output
rlabel metal2 s 18502 0 18530 82 6 output_thermometer_o[16]
port 128 nsew signal output
rlabel metal2 s 18778 41670 18806 42000 6 output_thermometer_o[158]
port 129 nsew signal output
rlabel metal2 s 18778 0 18806 218 6 output_thermometer_o[45]
port 130 nsew signal output
rlabel metal2 s 19054 41670 19082 42000 6 output_thermometer_o[87]
port 131 nsew signal output
rlabel metal2 s 19054 0 19082 82 6 output_thermometer_o[149]
port 132 nsew signal output
rlabel metal2 s 19330 41744 19358 42000 6 output_thermometer_o[237]
port 133 nsew signal output
rlabel metal2 s 19330 0 19358 144 6 output_thermometer_o[224]
port 134 nsew signal output
rlabel metal2 s 19606 41670 19634 42000 6 output_thermometer_o[154]
port 135 nsew signal output
rlabel metal2 s 19606 0 19634 82 6 output_thermometer_o[98]
port 136 nsew signal output
rlabel metal2 s 19882 41670 19910 42000 6 output_thermometer_o[19]
port 137 nsew signal output
rlabel metal2 s 19882 0 19910 82 6 output_thermometer_o[222]
port 138 nsew signal output
rlabel metal2 s 20158 41670 20186 42000 6 output_thermometer_o[181]
port 139 nsew signal output
rlabel metal2 s 20158 0 20186 82 6 output_thermometer_o[35]
port 140 nsew signal output
rlabel metal2 s 20434 41670 20462 42000 6 output_thermometer_o[207]
port 141 nsew signal output
rlabel metal2 s 20434 0 20462 82 6 output_thermometer_o[124]
port 142 nsew signal output
rlabel metal2 s 20710 41670 20738 42000 6 output_thermometer_o[140]
port 143 nsew signal output
rlabel metal2 s 20710 0 20738 218 6 output_thermometer_o[25]
port 144 nsew signal output
rlabel metal2 s 20986 41670 21014 42000 6 output_thermometer_o[126]
port 145 nsew signal output
rlabel metal2 s 20986 0 21014 218 6 output_thermometer_o[68]
port 146 nsew signal output
rlabel metal2 s 21262 41806 21290 42000 6 output_thermometer_o[143]
port 147 nsew signal output
rlabel metal2 s 21262 0 21290 82 6 output_thermometer_o[175]
port 148 nsew signal output
rlabel metal2 s 21538 41670 21566 42000 6 output_thermometer_o[13]
port 149 nsew signal output
rlabel metal2 s 21538 0 21566 82 6 output_thermometer_o[178]
port 150 nsew signal output
rlabel metal2 s 21814 41806 21842 42000 6 output_thermometer_o[248]
port 151 nsew signal output
rlabel metal2 s 21814 0 21842 218 6 output_thermometer_o[131]
port 152 nsew signal output
rlabel metal2 s 22090 41670 22118 42000 6 output_thermometer_o[95]
port 153 nsew signal output
rlabel metal2 s 22090 0 22118 218 6 output_thermometer_o[156]
port 154 nsew signal output
rlabel metal2 s 22366 41670 22394 42000 6 output_thermometer_o[89]
port 155 nsew signal output
rlabel metal2 s 22366 0 22394 218 6 output_thermometer_o[176]
port 156 nsew signal output
rlabel metal2 s 22642 41670 22670 42000 6 output_thermometer_o[205]
port 157 nsew signal output
rlabel metal2 s 22642 0 22670 82 6 output_thermometer_o[62]
port 158 nsew signal output
rlabel metal2 s 22918 41670 22946 42000 6 output_thermometer_o[39]
port 159 nsew signal output
rlabel metal2 s 22918 0 22946 82 6 output_thermometer_o[99]
port 160 nsew signal output
rlabel metal2 s 23194 41670 23222 42000 6 output_thermometer_o[41]
port 161 nsew signal output
rlabel metal2 s 23194 0 23222 82 6 output_thermometer_o[104]
port 162 nsew signal output
rlabel metal2 s 23470 41670 23498 42000 6 output_thermometer_o[169]
port 163 nsew signal output
rlabel metal2 s 23470 0 23498 82 6 output_binary_o[0]
port 164 nsew signal output
rlabel metal2 s 23746 41670 23774 42000 6 output_thermometer_o[186]
port 165 nsew signal output
rlabel metal2 s 23746 0 23774 218 6 output_thermometer_o[180]
port 166 nsew signal output
rlabel metal2 s 24022 41670 24050 42000 6 output_thermometer_o[214]
port 167 nsew signal output
rlabel metal2 s 24022 0 24050 82 6 output_thermometer_o[63]
port 168 nsew signal output
rlabel metal2 s 24298 41670 24326 42000 6 output_thermometer_o[206]
port 169 nsew signal output
rlabel metal2 s 24298 0 24326 82 6 output_thermometer_o[128]
port 170 nsew signal output
rlabel metal2 s 24574 41670 24602 42000 6 output_thermometer_o[228]
port 171 nsew signal output
rlabel metal2 s 24574 0 24602 218 6 output_thermometer_o[55]
port 172 nsew signal output
rlabel metal2 s 24850 41670 24878 42000 6 output_thermometer_o[220]
port 173 nsew signal output
rlabel metal2 s 24850 0 24878 218 6 output_thermometer_o[111]
port 174 nsew signal output
rlabel metal2 s 25126 41670 25154 42000 6 output_thermometer_o[247]
port 175 nsew signal output
rlabel metal2 s 25126 0 25154 218 6 output_thermometer_o[183]
port 176 nsew signal output
rlabel metal2 s 25402 41670 25430 42000 6 output_thermometer_o[219]
port 177 nsew signal output
rlabel metal2 s 25402 0 25430 218 6 output_thermometer_o[58]
port 178 nsew signal output
rlabel metal2 s 25678 41670 25706 42000 6 output_thermometer_o[114]
port 179 nsew signal output
rlabel metal2 s 25678 0 25706 212 6 output_thermometer_o[252]
port 180 nsew signal output
rlabel metal2 s 25954 41670 25982 42000 6 output_thermometer_o[167]
port 181 nsew signal output
rlabel metal2 s 25954 0 25982 252 6 output_thermometer_o[49]
port 182 nsew signal output
rlabel metal2 s 26230 41670 26258 42000 6 output_thermometer_o[159]
port 183 nsew signal output
rlabel metal2 s 26230 0 26258 82 6 output_thermometer_o[120]
port 184 nsew signal output
rlabel metal2 s 26506 41670 26534 42000 6 output_thermometer_o[78]
port 185 nsew signal output
rlabel metal2 s 26506 0 26534 218 6 output_thermometer_o[152]
port 186 nsew signal output
rlabel metal2 s 26782 41670 26810 42000 6 output_thermometer_o[189]
port 187 nsew signal output
rlabel metal2 s 26782 0 26810 218 6 output_thermometer_o[103]
port 188 nsew signal output
rlabel metal2 s 27058 41670 27086 42000 6 output_thermometer_o[106]
port 189 nsew signal output
rlabel metal2 s 27058 0 27086 82 6 output_thermometer_o[233]
port 190 nsew signal output
rlabel metal2 s 27334 41670 27362 42000 6 output_thermometer_o[155]
port 191 nsew signal output
rlabel metal2 s 27334 0 27362 218 6 output_thermometer_o[34]
port 192 nsew signal output
rlabel metal2 s 27610 41670 27638 42000 6 output_thermometer_o[138]
port 193 nsew signal output
rlabel metal2 s 27610 0 27638 82 6 output_thermometer_o[48]
port 194 nsew signal output
rlabel metal2 s 27886 41670 27914 42000 6 output_binary_o[1]
port 195 nsew signal output
rlabel metal2 s 27886 0 27914 82 6 output_thermometer_o[225]
port 196 nsew signal output
rlabel metal2 s 28162 41670 28190 42000 6 output_thermometer_o[121]
port 197 nsew signal output
rlabel metal2 s 28162 0 28190 218 6 output_thermometer_o[10]
port 198 nsew signal output
rlabel metal2 s 28438 41670 28466 42000 6 output_thermometer_o[77]
port 199 nsew signal output
rlabel metal2 s 28438 0 28466 82 6 output_thermometer_o[170]
port 200 nsew signal output
rlabel metal2 s 28714 41670 28742 42000 6 output_thermometer_o[141]
port 201 nsew signal output
rlabel metal2 s 28714 0 28742 82 6 output_thermometer_o[40]
port 202 nsew signal output
rlabel metal2 s 28990 41670 29018 42000 6 output_thermometer_o[216]
port 203 nsew signal output
rlabel metal2 s 28990 0 29018 82 6 output_thermometer_o[139]
port 204 nsew signal output
rlabel metal2 s 29266 41670 29294 42000 6 output_thermometer_o[210]
port 205 nsew signal output
rlabel metal2 s 29266 0 29294 82 6 output_thermometer_o[42]
port 206 nsew signal output
rlabel metal2 s 29542 41670 29570 42000 6 output_thermometer_o[150]
port 207 nsew signal output
rlabel metal2 s 29542 0 29570 252 6 output_thermometer_o[88]
port 208 nsew signal output
rlabel metal2 s 29818 41744 29846 42000 6 output_thermometer_o[240]
port 209 nsew signal output
rlabel metal2 s 29818 0 29846 82 6 output_thermometer_o[1]
port 210 nsew signal output
rlabel metal2 s 30094 41670 30122 42000 6 output_thermometer_o[66]
port 211 nsew signal output
rlabel metal2 s 30094 0 30122 218 6 output_thermometer_o[36]
port 212 nsew signal output
rlabel metal2 s 30370 41670 30398 42000 6 output_thermometer_o[127]
port 213 nsew signal output
rlabel metal2 s 30370 0 30398 82 6 output_thermometer_o[177]
port 214 nsew signal output
rlabel metal2 s 30646 41670 30674 42000 6 output_thermometer_o[148]
port 215 nsew signal output
rlabel metal2 s 30646 0 30674 82 6 output_thermometer_o[239]
port 216 nsew signal output
rlabel metal2 s 30922 41670 30950 42000 6 output_thermometer_o[255]
port 217 nsew signal output
rlabel metal2 s 30922 0 30950 82 6 output_thermometer_o[71]
port 218 nsew signal output
rlabel metal2 s 31198 41670 31226 42000 6 output_thermometer_o[133]
port 219 nsew signal output
rlabel metal2 s 31198 0 31226 82 6 output_thermometer_o[91]
port 220 nsew signal output
rlabel metal2 s 31474 41670 31502 42000 6 output_thermometer_o[22]
port 221 nsew signal output
rlabel metal2 s 31474 0 31502 218 6 output_thermometer_o[65]
port 222 nsew signal output
rlabel metal2 s 31750 41880 31778 42000 6 output_thermometer_o[75]
port 223 nsew signal output
rlabel metal2 s 31750 0 31778 82 6 output_thermometer_o[192]
port 224 nsew signal output
rlabel metal2 s 32026 41670 32054 42000 6 output_thermometer_o[51]
port 225 nsew signal output
rlabel metal2 s 32026 0 32054 218 6 output_thermometer_o[171]
port 226 nsew signal output
rlabel metal2 s 32302 41670 32330 42000 6 output_thermometer_o[254]
port 227 nsew signal output
rlabel metal2 s 32302 0 32330 82 6 output_thermometer_o[28]
port 228 nsew signal output
rlabel metal2 s 32578 41670 32606 42000 6 output_thermometer_o[122]
port 229 nsew signal output
rlabel metal2 s 32578 0 32606 82 6 output_thermometer_o[70]
port 230 nsew signal output
rlabel metal2 s 32854 41670 32882 42000 6 output_thermometer_o[46]
port 231 nsew signal output
rlabel metal2 s 32854 0 32882 218 6 output_thermometer_o[100]
port 232 nsew signal output
rlabel metal2 s 33130 41744 33158 42000 6 output_thermometer_o[56]
port 233 nsew signal output
rlabel metal2 s 33130 0 33158 212 6 output_thermometer_o[172]
port 234 nsew signal output
rlabel metal2 s 33406 41806 33434 42000 6 output_thermometer_o[135]
port 235 nsew signal output
rlabel metal2 s 33406 0 33434 82 6 output_thermometer_o[184]
port 236 nsew signal output
rlabel metal2 s 33682 41812 33710 42000 6 output_thermometer_o[173]
port 237 nsew signal output
rlabel metal2 s 33682 0 33710 82 6 output_thermometer_o[85]
port 238 nsew signal output
rlabel metal2 s 33958 41670 33986 42000 6 output_thermometer_o[38]
port 239 nsew signal output
rlabel metal2 s 33958 0 33986 218 6 output_thermometer_o[52]
port 240 nsew signal output
rlabel metal2 s 34234 41670 34262 42000 6 output_thermometer_o[238]
port 241 nsew signal output
rlabel metal2 s 34234 0 34262 82 6 output_thermometer_o[92]
port 242 nsew signal output
rlabel metal2 s 34510 41670 34538 42000 6 output_thermometer_o[165]
port 243 nsew signal output
rlabel metal2 s 34510 0 34538 82 6 output_thermometer_o[223]
port 244 nsew signal output
rlabel metal2 s 34786 41670 34814 42000 6 output_thermometer_o[246]
port 245 nsew signal output
rlabel metal2 s 34786 0 34814 218 6 output_thermometer_o[118]
port 246 nsew signal output
rlabel metal2 s 35062 41670 35090 42000 6 output_thermometer_o[50]
port 247 nsew signal output
rlabel metal2 s 35062 0 35090 82 6 output_thermometer_o[202]
port 248 nsew signal output
rlabel metal2 s 35338 41806 35366 42000 6 output_thermometer_o[113]
port 249 nsew signal output
rlabel metal2 s 35338 0 35366 218 6 output_thermometer_o[80]
port 250 nsew signal output
rlabel metal2 s 35614 41670 35642 42000 6 output_thermometer_o[231]
port 251 nsew signal output
rlabel metal2 s 35614 0 35642 218 6 output_thermometer_o[153]
port 252 nsew signal output
rlabel metal2 s 35890 41670 35918 42000 6 output_thermometer_o[203]
port 253 nsew signal output
rlabel metal2 s 35890 0 35918 82 6 output_thermometer_o[6]
port 254 nsew signal output
rlabel metal2 s 36166 41670 36194 42000 6 output_thermometer_o[44]
port 255 nsew signal output
rlabel metal2 s 36166 0 36194 218 6 output_thermometer_o[0]
port 256 nsew signal output
rlabel metal2 s 36442 41744 36470 42000 6 output_thermometer_o[108]
port 257 nsew signal output
rlabel metal2 s 36442 0 36470 218 6 output_thermometer_o[24]
port 258 nsew signal output
rlabel metal2 s 36718 41670 36746 42000 6 en_o
port 259 nsew signal output
rlabel metal3 s 79760 19036 80000 19156 6 clk_i
port 260 nsew signal input
rlabel metal3 s 79760 19308 80000 19428 6 rst_ni
port 261 nsew signal input
rlabel metal3 s 79760 19580 80000 19700 6 randomise_en_i
port 262 nsew signal input
rlabel metal3 s 79760 19852 80000 19972 6 en_i
port 263 nsew signal input
rlabel metal3 s 79760 20124 80000 20244 6 input_binary_i[0]
port 264 nsew signal input
rlabel metal3 s 79760 20396 80000 20516 6 input_binary_i[1]
port 265 nsew signal input
rlabel metal3 s 79760 20668 80000 20788 6 input_binary_i[2]
port 266 nsew signal input
rlabel metal3 s 79760 20940 80000 21060 6 input_binary_i[3]
port 267 nsew signal input
rlabel metal3 s 79760 21212 80000 21332 6 input_binary_i[4]
port 268 nsew signal input
rlabel metal3 s 79760 21484 80000 21604 6 input_binary_i[5]
port 269 nsew signal input
rlabel metal3 s 79760 21756 80000 21876 6 input_binary_i[6]
port 270 nsew signal input
rlabel metal3 s 79760 22028 80000 22148 6 input_binary_i[7]
port 271 nsew signal input
rlabel metal3 s 79760 22300 80000 22420 6 input_binary_i[8]
port 272 nsew signal input
rlabel metal3 s 79760 22572 80000 22692 6 input_binary_i[9]
port 273 nsew signal input
rlabel metal4 s 65648 2128 65968 39760 6 VPWR
port 274 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 39760 6 VPWR
port 275 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 39760 6 VPWR
port 276 nsew power bidirectional
rlabel metal5 s 1104 35934 78844 36254 6 VPWR
port 277 nsew power bidirectional
rlabel metal5 s 1104 5298 78844 5618 6 VPWR
port 278 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 39760 6 VGND
port 279 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 39760 6 VGND
port 280 nsew ground bidirectional
rlabel metal5 s 1104 20616 78844 20936 6 VGND
port 281 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 80000 42000
string LEFview TRUE
string GDS_FILE /amsat_txrx_ic/design/dac_digital_interface/runs/16-05_11-04/results/magic/dac_digital_interface.gds
string GDS_END 8231378
string GDS_START 507552
<< end >>

