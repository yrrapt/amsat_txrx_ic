**.subckt bandgap_core_stability_ptat
x1 net4 ptat net13 net14 net17 GND bandgap_opamp
x2 net4 ctat net5 net1 net7 GND bandgap_opamp
XM3 net6 net6 GND GND sky130_fd_pr__nfet_01v8_lvt W=7 L=8 ad=2.03 pd=14.58 as=2.03 ps=14.58
+ nrd=0.041428571428571426 nrs=0.041428571428571426 sa=0 sb=0 sd=0 nf=1 mult=2 m=2
XM1 cas net6 GND GND sky130_fd_pr__nfet_01v8_lvt W=7 L=8 ad=2.03 pd=14.58 as=2.03 ps=14.58
+ nrd=0.041428571428571426 nrs=0.041428571428571426 sa=0 sb=0 sd=0 nf=1 mult=2 m=2
.save v( net2 )
.save v( net1 )
.save v( net5 )
.save v( cas )
v2 net11 net17 0
x5 net4 ptat cas net8 bandgap_cascurr_cell m=8
x6 net4 ptat cas net9 bandgap_cascurr_cell m=8
x7 net4 ctat cas net10 bandgap_cascurr_cell m=8
x10 net4 ptat cas net6 bandgap_cascurr_cell m=2
x11 net4 ctat cas net6 bandgap_cascurr_cell m=2
XQ1 GND GND net3 GND sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8
XQ2 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
v3 net8 net2 0
v5 net9 net1 0
v6 net10 net5 0
C1 ctat net1 1m m=1
XR1 net3 net2 GND sky130_fd_pr__res_xhigh_po W=1 L=3.25 m=1
XR2 GND net5 GND sky130_fd_pr__res_xhigh_po W=1 L=28.6 m=1
.save v( net11 )
.save v( ctat )
x8 net4 net4 bmr_biasv GND bandgap_bmr
XMcurr net11 bmr_biasv net4 net4 sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr1 net7 bmr_biasv net4 net4 sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
Vdd net4 GND {vdd} 
Vin net12 GND dc=0 ac=1
XMcurr2 net4 ptat net4 net4 sky130_fd_pr__pfet_01v8_lvt W=7 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
Vin1 net15 GND dc=0 ac=-1
E1 ac GND net2 net1 1
Vctl4 ctl_ptat[4] GND {ctl4} 
Vctl3 ctl_ptat[3] GND {ctl3} 
Vctl2 ctl_ptat[2] GND {ctl2} 
Vctl1 ctl_ptat[1] GND {ctl1} 
Vctl0 ctl_ptat[0] GND {ctl0} 
R3 net2 net13 1u m=1 ac=1G
R5 net1 net14 1u m=1 ac=1G
R4 net12 net13 1G m=1 ac=1u
R6 net15 net14 1G m=1 ac=1u
XM8 net16 cas net4 net4 sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMcpdiff1 cas cas net16 net4 sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
**** begin user architecture code


.temp 27

.lib sky130_fd_pr/models/sky130.lib.spice tt
.include sky130_fd_pr/models/sky130_fd_pr__model__pnp.model.spice

.param vdd=1.8

.param ctl4=0
.param ctl3=0
.param ctl2=0
.param ctl1=0
.param ctl0=0

.save all

*.op
.ac dec 10 1 1G

*.control
*   run
*   setplot ac1
*   set units=degrees
*   gnuplot bandgap_core_stability2 db(fb) ph(fb)
*.endc


**** end user architecture code
**.ends

* expanding   symbol:  bandgap_opamp/bandgap_opamp.sym # of pins=6

.subckt bandgap_opamp  vdd out inp inn bias gnd
*.ipin inp
*.ipin inn
*.ipin bias
*.opin out
*.iopin vdd
*.iopin gnd
XMmpdiff net9 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=32 m=32 
XMmpr net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMmnr bias bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=2 m=2
XMmnb net2 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=2 m=2
XMtrioden net11 net5 gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=8 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=1 m=1
XMmpa net10 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcpdiff net1 net8 net9 vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=32 m=32 
XMmna net8 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=2 m=2
XMtriodep net12 net8 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMcpa net5 net8 net10 vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcasba net5 net5 net11 gnd sky130_fd_pr__nfet_01v8_lvt W=5 L=4 ad=1.45 pd=10.58 as=1.45 ps=10.58
+ nrd=0.057999999999999996 nrs=0.057999999999999996 sa=0 sb=0 sd=0 nf=1 mult=8 m=8
.save v( net3 )
XMcasn net7 net5 net4 gnd sky130_fd_pr__nfet_01v8_lvt W=5 L=4 ad=1.45 pd=10.58 as=1.45 ps=10.58
+ nrd=0.057999999999999996 nrs=0.057999999999999996 sa=0 sb=0 sd=0 nf=1 mult=8 m=8
XMcasp net6 net5 net3 gnd sky130_fd_pr__nfet_01v8_lvt W=5 L=4 ad=1.45 pd=10.58 as=1.45 ps=10.58
+ nrd=0.057999999999999996 nrs=0.057999999999999996 sa=0 sb=0 sd=0 nf=1 mult=8 m=8
XMloadmp net13 net6 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMloadmn net14 net6 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMloadcn net7 net8 net14 vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=10 m=10 
XMloadcp net6 net8 net13 vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=10 m=10 
XMmfn net4 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=8 m=8
XMmfp net3 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ nrd=0.145 nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=8 m=8
XMdiffn net4 inp net1 net1 sky130_fd_pr__pfet_01v8_lvt W=7 L=0.35 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=64 m=64 
XMdiffp net3 inn net1 net1 sky130_fd_pr__pfet_01v8_lvt W=7 L=0.35 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=64 m=64 
.save v( net5 )
.save v( net1 )
.save v( net8 )
.save v( net2 )
.save v( net14 )
.save v( net6 )
XMcpdiff1 net8 net8 net12 vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
.save v( net4 )
XMmnc out bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad=0.58 pd=4.58 as=0.58 ps=4.58 nrd=0.145
+ nrs=0.145 sa=0 sb=0 sd=0 nf=1 mult=32 m=32
XMgain out net7 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XC1 out out sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1
.ends


* expanding   symbol:  bandgap_cascurr_cell/bandgap_cascurr_cell.sym # of pins=4

.subckt bandgap_cascurr_cell  vdd curr cas out
*.iopin vdd
*.ipin curr
*.ipin cas
*.opin out
XMcurr net1 curr vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMcas out cas net1 vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
.save v( net1 )
.ends


* expanding   symbol:  bandgap_bmr/bandgap_bmr.sym # of pins=4

.subckt bandgap_bmr  vdd en biasv vss
*.iopin vdd
*.iopin vss
*.opin biasv
*.ipin en
XMdiff_n2 biasv net1 net2 vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XR1 vss net2 vss sky130_fd_pr__res_xhigh_po W=1 L=5 m=1
XMdiff_n1 net1 net1 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_p2 biasv biasv vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_p1 net1 biasv vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMsw_start biasv net3 net1 vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMdiff_n3 net3 net1 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_bias net3 net3 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en2 biasv en vdd vdd sky130_fd_pr__pfet_01v8_lvt W=0.42 L=0.35 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en1 net3 en vdd vdd sky130_fd_pr__pfet_01v8_lvt W=0.42 L=0.35 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XCcomp biasv net1 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1
XMdum vss net1 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=5 m=5 
XCfilt biasv vdd sky130_fd_pr__cap_mim_m3_1 W=7.7 L=7.2 MF=1
.ends

.GLOBAL GND
.end
