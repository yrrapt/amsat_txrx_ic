* NGSPICE file created from dac_digital_interface.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

.subckt dac_digital_interface output_binary_o[0] output_binary_o[1] output_thermometer_o[252]
+ output_thermometer_o[29] output_thermometer_o[58] output_thermometer_o[91] output_thermometer_o[64]
+ output_thermometer_o[15] output_thermometer_o[28] output_thermometer_o[19] output_thermometer_o[128]
+ output_thermometer_o[145] output_thermometer_o[43] output_thermometer_o[239] output_thermometer_o[68]
+ output_thermometer_o[164] output_thermometer_o[131] output_thermometer_o[72] output_thermometer_o[99]
+ output_thermometer_o[143] output_thermometer_o[193] output_thermometer_o[229] output_thermometer_o[67]
+ output_thermometer_o[176] output_thermometer_o[125] output_thermometer_o[59] output_thermometer_o[202]
+ output_thermometer_o[78] output_thermometer_o[116] output_thermometer_o[21] output_thermometer_o[41]
+ output_thermometer_o[3] output_thermometer_o[39] output_thermometer_o[18] output_thermometer_o[77]
+ output_thermometer_o[249] output_thermometer_o[34] output_thermometer_o[102] output_thermometer_o[124]
+ output_thermometer_o[106] output_thermometer_o[14] output_thermometer_o[217] output_thermometer_o[112]
+ output_thermometer_o[156] output_thermometer_o[189] output_thermometer_o[196] output_thermometer_o[152]
+ output_thermometer_o[215] output_thermometer_o[92] output_thermometer_o[171] output_thermometer_o[94]
+ output_thermometer_o[42] output_thermometer_o[79] output_thermometer_o[144] output_thermometer_o[150]
+ output_thermometer_o[137] output_thermometer_o[83] output_thermometer_o[245] output_thermometer_o[82]
+ output_thermometer_o[180] output_thermometer_o[54] output_thermometer_o[123] output_thermometer_o[37]
+ output_thermometer_o[26] output_thermometer_o[46] output_thermometer_o[11] output_thermometer_o[88]
+ output_thermometer_o[121] output_thermometer_o[186] output_thermometer_o[212] output_thermometer_o[194]
+ output_thermometer_o[244] output_thermometer_o[182] output_thermometer_o[120] output_thermometer_o[52]
+ output_thermometer_o[223] output_thermometer_o[25] output_thermometer_o[172] output_thermometer_o[197]
+ output_thermometer_o[232] output_thermometer_o[242] output_thermometer_o[203] output_thermometer_o[95]
+ output_thermometer_o[130] output_thermometer_o[195] output_thermometer_o[228] output_thermometer_o[230]
+ output_thermometer_o[63] output_thermometer_o[9] output_thermometer_o[201] output_thermometer_o[183]
+ output_thermometer_o[237] output_thermometer_o[44] output_thermometer_o[134] output_thermometer_o[35]
+ output_thermometer_o[113] output_thermometer_o[73] output_thermometer_o[4] output_thermometer_o[219]
+ output_thermometer_o[0] output_thermometer_o[221] output_thermometer_o[96] output_thermometer_o[74]
+ output_thermometer_o[207] output_thermometer_o[127] output_thermometer_o[20] output_thermometer_o[24]
+ output_thermometer_o[246] output_thermometer_o[153] output_thermometer_o[154] output_thermometer_o[155]
+ output_thermometer_o[170] output_thermometer_o[160] output_thermometer_o[100] output_thermometer_o[85]
+ output_thermometer_o[192] output_thermometer_o[48] output_thermometer_o[139] output_thermometer_o[248]
+ output_thermometer_o[190] output_thermometer_o[109] output_thermometer_o[81] output_thermometer_o[12]
+ output_thermometer_o[133] output_thermometer_o[167] output_thermometer_o[204] output_thermometer_o[222]
+ output_thermometer_o[142] output_thermometer_o[199] output_thermometer_o[240] output_thermometer_o[103]
+ output_thermometer_o[138] output_thermometer_o[97] output_thermometer_o[89] output_thermometer_o[175]
+ output_thermometer_o[84] output_thermometer_o[250] output_thermometer_o[251] output_thermometer_o[162]
+ output_thermometer_o[10] output_thermometer_o[6] output_thermometer_o[148] output_thermometer_o[110]
+ output_thermometer_o[98] output_thermometer_o[146] output_thermometer_o[225] output_thermometer_o[108]
+ output_thermometer_o[53] output_thermometer_o[115] output_thermometer_o[62] output_thermometer_o[169]
+ output_thermometer_o[5] output_thermometer_o[140] output_thermometer_o[49] output_thermometer_o[149]
+ output_thermometer_o[118] output_thermometer_o[191] output_thermometer_o[168] output_thermometer_o[135]
+ output_thermometer_o[141] output_thermometer_o[90] output_thermometer_o[2] output_thermometer_o[213]
+ output_thermometer_o[93] output_thermometer_o[173] output_thermometer_o[55] output_thermometer_o[105]
+ output_thermometer_o[101] output_thermometer_o[111] output_thermometer_o[205] output_thermometer_o[132]
+ output_thermometer_o[159] output_thermometer_o[32] output_thermometer_o[233] output_thermometer_o[208]
+ output_thermometer_o[16] output_thermometer_o[163] output_thermometer_o[178] output_thermometer_o[86]
+ output_thermometer_o[188] output_thermometer_o[200] output_thermometer_o[104] output_thermometer_o[136]
+ output_thermometer_o[33] output_thermometer_o[174] output_thermometer_o[209] output_thermometer_o[206]
+ output_thermometer_o[129] output_thermometer_o[70] output_thermometer_o[38] output_thermometer_o[187]
+ output_thermometer_o[23] output_thermometer_o[224] output_thermometer_o[179] output_thermometer_o[117]
+ output_thermometer_o[236] output_thermometer_o[114] output_thermometer_o[13] output_thermometer_o[177]
+ output_thermometer_o[231] output_thermometer_o[45] output_thermometer_o[254] output_thermometer_o[161]
+ output_thermometer_o[238] output_thermometer_o[47] output_thermometer_o[147] output_thermometer_o[30]
+ output_thermometer_o[218] output_thermometer_o[211] output_thermometer_o[40] output_thermometer_o[57]
+ output_thermometer_o[8] output_thermometer_o[50] output_thermometer_o[36] output_thermometer_o[210]
+ output_thermometer_o[27] output_thermometer_o[51] output_thermometer_o[165] output_thermometer_o[60]
+ output_thermometer_o[65] output_thermometer_o[253] output_thermometer_o[71] output_thermometer_o[181]
+ output_thermometer_o[107] output_thermometer_o[234] output_thermometer_o[17] output_thermometer_o[216]
+ output_thermometer_o[56] output_thermometer_o[119] output_thermometer_o[166] output_thermometer_o[61]
+ output_thermometer_o[126] output_thermometer_o[185] output_thermometer_o[241] output_thermometer_o[220]
+ output_thermometer_o[243] output_thermometer_o[87] output_thermometer_o[122] output_thermometer_o[1]
+ output_thermometer_o[151] output_thermometer_o[76] output_thermometer_o[22] output_thermometer_o[66]
+ output_thermometer_o[158] output_thermometer_o[198] output_thermometer_o[31] output_thermometer_o[184]
+ output_thermometer_o[80] output_thermometer_o[7] output_thermometer_o[75] output_thermometer_o[247]
+ output_thermometer_o[157] output_thermometer_o[226] output_thermometer_o[227] output_thermometer_o[69]
+ output_thermometer_o[255] output_thermometer_o[214] output_thermometer_o[235] clk_i
+ rst_ni randomise_en_i input_binary_i[0] input_binary_i[1] input_binary_i[2] input_binary_i[3]
+ input_binary_i[4] input_binary_i[5] input_binary_i[6] input_binary_i[7] input_binary_i[8]
+ input_binary_i[9] VPWR VGND
X_3155_ _2687_/Y _2685_/Y _3347_/S VGND VGND VPWR VPWR _3155_/X sky130_fd_sc_hd__mux2_4
XFILLER_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2106_ _1777_/X _2790_/B _2097_/X _3021_/A _2105_/X VGND VGND VPWR VPWR _2106_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_54_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3086_ _3110_/A VGND VGND VPWR VPWR _3107_/A sky130_fd_sc_hd__clkbuf_2
X_2037_ _1992_/X _2019_/X _2020_/X _2526_/A _2023_/X VGND VGND VPWR VPWR _3000_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_54_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2939_ _2939_/A VGND VGND VPWR VPWR _3001_/A sky130_fd_sc_hd__buf_2
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2724_ _2724_/A _2956_/B VGND VGND VPWR VPWR _2724_/X sky130_fd_sc_hd__or2_1
X_2655_ _3111_/B _2653_/X _2171_/A _2881_/B _2654_/X VGND VGND VPWR VPWR _2655_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1606_ _2401_/A _2407_/A VGND VGND VPWR VPWR _2669_/B sky130_fd_sc_hd__nor2_2
X_2586_ _3027_/A VGND VGND VPWR VPWR _2662_/A sky130_fd_sc_hd__clkbuf_2
X_3207_ _2876_/Y _2335_/A _3351_/S VGND VGND VPWR VPWR _3207_/X sky130_fd_sc_hd__mux2_2
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3138_ _2628_/Y _2625_/Y _3330_/S VGND VGND VPWR VPWR _3138_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3069_ _3108_/A _3069_/B VGND VGND VPWR VPWR _3069_/X sky130_fd_sc_hd__or2_1
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2440_ _2440_/A _2803_/B VGND VGND VPWR VPWR _2440_/X sky130_fd_sc_hd__or2_1
X_2371_ _2380_/A _2373_/A VGND VGND VPWR VPWR _2656_/B sky130_fd_sc_hd__nor2_4
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2707_ _2718_/A _2707_/B VGND VGND VPWR VPWR _2707_/Y sky130_fd_sc_hd__nor2_1
Xoutput253 _3204_/X VGND VGND VPWR VPWR output_thermometer_o[76] sky130_fd_sc_hd__clkbuf_2
Xoutput231 _3188_/X VGND VGND VPWR VPWR output_thermometer_o[60] sky130_fd_sc_hd__clkbuf_2
Xoutput220 _3346_/X VGND VGND VPWR VPWR output_thermometer_o[218] sky130_fd_sc_hd__clkbuf_2
X_2638_ _3093_/B _2630_/X _2626_/X _2868_/B _2637_/X VGND VGND VPWR VPWR _2638_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput242 _3294_/X VGND VGND VPWR VPWR output_thermometer_o[166] sky130_fd_sc_hd__clkbuf_2
X_2569_ _2811_/B _2390_/X _3042_/B _2206_/X VGND VGND VPWR VPWR _2569_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput264 _3285_/X VGND VGND VPWR VPWR output_thermometer_o[157] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1940_ _1964_/A _1940_/B VGND VGND VPWR VPWR _2737_/B sky130_fd_sc_hd__nor2_2
X_1871_ _2157_/A VGND VGND VPWR VPWR _1871_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2423_ _2422_/X _2916_/B _2917_/A _2415_/X VGND VGND VPWR VPWR _2423_/X sky130_fd_sc_hd__o22a_1
X_2354_ _2291_/X _2650_/A _2898_/A VGND VGND VPWR VPWR _2878_/B sky130_fd_sc_hd__o21a_1
X_2285_ _2286_/A _2317_/B VGND VGND VPWR VPWR _3083_/B sky130_fd_sc_hd__nor2_2
XFILLER_37_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2070_ _2081_/A _2070_/B VGND VGND VPWR VPWR _2781_/B sky130_fd_sc_hd__nor2_4
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2972_ _2975_/A _2972_/B VGND VGND VPWR VPWR _2972_/X sky130_fd_sc_hd__or2_1
X_1923_ _1871_/X _2486_/A _1875_/X VGND VGND VPWR VPWR _1927_/B sky130_fd_sc_hd__o21ai_2
X_1854_ _2087_/A VGND VGND VPWR VPWR _1854_/X sky130_fd_sc_hd__buf_2
X_1785_ _2391_/A VGND VGND VPWR VPWR _2301_/A sky130_fd_sc_hd__clkbuf_2
X_2406_ _2406_/A VGND VGND VPWR VPWR _2406_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3386_ _3408_/CLK input7/X VGND VGND VPWR VPWR _3386_/Q sky130_fd_sc_hd__dfxtp_1
X_2337_ _2324_/X _2327_/Y _2336_/X VGND VGND VPWR VPWR _2337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2268_ _2329_/B _2268_/B VGND VGND VPWR VPWR _2269_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2199_ _2219_/A _2199_/B VGND VGND VPWR VPWR _3054_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 _3295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ _1570_/A _2329_/B VGND VGND VPWR VPWR _1601_/A sky130_fd_sc_hd__or2_1
X_3240_ _2995_/Y _2992_/Y _3370_/S VGND VGND VPWR VPWR _3240_/X sky130_fd_sc_hd__mux2_2
X_3171_ _2745_/Y _2741_/Y _3365_/S VGND VGND VPWR VPWR _3171_/X sky130_fd_sc_hd__mux2_4
XFILLER_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2122_ _2156_/A _2122_/B VGND VGND VPWR VPWR _2798_/B sky130_fd_sc_hd__nor2_4
XFILLER_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2053_ _2034_/X _3003_/B _2025_/X _2772_/B _2052_/X VGND VGND VPWR VPWR _2053_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2955_ _2967_/A _2955_/B VGND VGND VPWR VPWR _2955_/Y sky130_fd_sc_hd__nor2_1
X_1906_ _1854_/X _2958_/B _1902_/X _2726_/B _1905_/X VGND VGND VPWR VPWR _1906_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2886_ _2886_/A _2886_/B VGND VGND VPWR VPWR _2886_/Y sky130_fd_sc_hd__nor2_1
X_1837_ _1843_/B VGND VGND VPWR VPWR _1838_/B sky130_fd_sc_hd__inv_2
X_1768_ _2185_/A _1769_/C VGND VGND VPWR VPWR _2434_/A sky130_fd_sc_hd__or2_2
X_1699_ _3385_/Q _3384_/Q _1847_/A VGND VGND VPWR VPWR _1759_/B sky130_fd_sc_hd__a21oi_2
X_3369_ _2525_/Y _2522_/Y _3374_/S VGND VGND VPWR VPWR _3369_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput20 _3143_/X VGND VGND VPWR VPWR output_thermometer_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput31 _3227_/X VGND VGND VPWR VPWR output_thermometer_o[99] sky130_fd_sc_hd__clkbuf_2
Xoutput42 _3149_/X VGND VGND VPWR VPWR output_thermometer_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput53 _3142_/X VGND VGND VPWR VPWR output_thermometer_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput75 _3165_/X VGND VGND VPWR VPWR output_thermometer_o[37] sky130_fd_sc_hd__clkbuf_2
Xoutput64 _3170_/X VGND VGND VPWR VPWR output_thermometer_o[42] sky130_fd_sc_hd__clkbuf_2
Xoutput86 _3248_/X VGND VGND VPWR VPWR output_thermometer_o[120] sky130_fd_sc_hd__clkbuf_2
Xoutput97 _3323_/X VGND VGND VPWR VPWR output_thermometer_o[195] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2740_ _2759_/A VGND VGND VPWR VPWR _2756_/A sky130_fd_sc_hd__clkbuf_2
X_2671_ _2900_/B _2545_/X _2670_/X VGND VGND VPWR VPWR _2671_/Y sky130_fd_sc_hd__o21ai_1
X_1622_ _2832_/A VGND VGND VPWR VPWR _1622_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3223_ _2933_/Y _2931_/Y _3351_/S VGND VGND VPWR VPWR _3223_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3154_ _2684_/Y _2681_/Y _3346_/S VGND VGND VPWR VPWR _3154_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2105_ _2548_/A _2993_/B _2879_/C VGND VGND VPWR VPWR _2105_/X sky130_fd_sc_hd__or3_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3085_ _3078_/X _2856_/B _3079_/X _2625_/B _3084_/X VGND VGND VPWR VPWR _3085_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2036_ _2036_/A VGND VGND VPWR VPWR _2526_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2938_ _2948_/A _2938_/B VGND VGND VPWR VPWR _2938_/Y sky130_fd_sc_hd__nor2_1
X_2869_ _3094_/B _2932_/B VGND VGND VPWR VPWR _2869_/X sky130_fd_sc_hd__or2_1
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2723_ _2723_/A VGND VGND VPWR VPWR _2723_/X sky130_fd_sc_hd__clkbuf_2
X_2654_ _2654_/A _2660_/B VGND VGND VPWR VPWR _2654_/X sky130_fd_sc_hd__or2_1
X_1605_ _1631_/A _1605_/B VGND VGND VPWR VPWR _2407_/A sky130_fd_sc_hd__or2_1
X_2585_ _2324_/X _1792_/Y _2581_/X _2584_/X VGND VGND VPWR VPWR _2585_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3206_ _2874_/Y _2871_/Y _3340_/S VGND VGND VPWR VPWR _3206_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3137_ _2624_/Y _2621_/Y _3330_/S VGND VGND VPWR VPWR _3137_/X sky130_fd_sc_hd__mux2_2
X_3068_ _3083_/A _3068_/B VGND VGND VPWR VPWR _3068_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2019_ _2141_/C VGND VGND VPWR VPWR _2019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ _2347_/X _2049_/A _1648_/A VGND VGND VPWR VPWR _2373_/A sky130_fd_sc_hd__o21ai_2
XFILLER_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2706_ _1816_/B _2704_/X _2935_/B _2673_/X _2705_/X VGND VGND VPWR VPWR _2706_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput210 _3141_/X VGND VGND VPWR VPWR output_thermometer_o[13] sky130_fd_sc_hd__clkbuf_2
X_2637_ _3094_/B _2641_/B VGND VGND VPWR VPWR _2637_/X sky130_fd_sc_hd__or2_1
Xoutput221 _3339_/X VGND VGND VPWR VPWR output_thermometer_o[211] sky130_fd_sc_hd__clkbuf_2
Xoutput243 _3189_/X VGND VGND VPWR VPWR output_thermometer_o[61] sky130_fd_sc_hd__clkbuf_2
Xoutput232 _3193_/X VGND VGND VPWR VPWR output_thermometer_o[65] sky130_fd_sc_hd__clkbuf_2
Xoutput254 _3150_/X VGND VGND VPWR VPWR output_thermometer_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput265 _3354_/X VGND VGND VPWR VPWR output_thermometer_o[226] sky130_fd_sc_hd__clkbuf_2
X_2568_ _2568_/A _2812_/A VGND VGND VPWR VPWR _2568_/Y sky130_fd_sc_hd__nor2_1
X_2499_ _2499_/A _2509_/B VGND VGND VPWR VPWR _2980_/B sky130_fd_sc_hd__or2_1
XFILLER_59_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1870_ _1854_/X _2948_/B _1842_/X _2714_/B _1869_/X VGND VGND VPWR VPWR _1870_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2422_ _2478_/A VGND VGND VPWR VPWR _2422_/X sky130_fd_sc_hd__buf_2
X_2353_ _2380_/A _2355_/A VGND VGND VPWR VPWR _2649_/B sky130_fd_sc_hd__nor2_4
X_2284_ _2184_/X _3084_/B _2185_/X VGND VGND VPWR VPWR _2856_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1999_ _2514_/A _2082_/A _2071_/C VGND VGND VPWR VPWR _1999_/X sky130_fd_sc_hd__or3_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2971_ _2985_/A _2971_/B VGND VGND VPWR VPWR _2971_/Y sky130_fd_sc_hd__nor2_1
X_1922_ _1922_/A VGND VGND VPWR VPWR _2486_/A sky130_fd_sc_hd__inv_2
X_1853_ _2832_/A VGND VGND VPWR VPWR _2087_/A sky130_fd_sc_hd__buf_2
X_1784_ _1777_/X _2697_/B _1660_/X _2931_/B _1783_/X VGND VGND VPWR VPWR _1784_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2405_ _2351_/X _2666_/B _2404_/X VGND VGND VPWR VPWR _2405_/Y sky130_fd_sc_hd__o21ai_1
X_3385_ _3408_/CLK input6/X VGND VGND VPWR VPWR _3385_/Q sky130_fd_sc_hd__dfxtp_2
X_2336_ _2328_/X _3101_/A _2331_/X _2335_/Y VGND VGND VPWR VPWR _2336_/X sky130_fd_sc_hd__o22a_1
X_2267_ _3080_/A _2618_/A VGND VGND VPWR VPWR _2851_/B sky130_fd_sc_hd__nor2_1
X_2198_ _2207_/A _2338_/A VGND VGND VPWR VPWR _2199_/B sky130_fd_sc_hd__or2_2
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 _3274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3170_ _2739_/Y _2737_/Y _3383_/S VGND VGND VPWR VPWR _3170_/X sky130_fd_sc_hd__mux2_2
X_2121_ _2155_/A _3029_/B VGND VGND VPWR VPWR _2121_/Y sky130_fd_sc_hd__nor2_1
X_2052_ _2530_/A _2061_/B VGND VGND VPWR VPWR _2052_/X sky130_fd_sc_hd__or2_1
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2954_ _2940_/X _1878_/B _2941_/X _2718_/B _2953_/X VGND VGND VPWR VPWR _2954_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1905_ _1917_/A _2476_/A _1954_/C VGND VGND VPWR VPWR _1905_/X sky130_fd_sc_hd__or3_2
X_2885_ _2882_/X _2652_/B _2840_/X _3112_/B _2884_/X VGND VGND VPWR VPWR _2885_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1836_ _1806_/X _2452_/A _2093_/A VGND VGND VPWR VPWR _1843_/B sky130_fd_sc_hd__o21ai_2
X_1767_ _2239_/A _1763_/B _1709_/X VGND VGND VPWR VPWR _1769_/C sky130_fd_sc_hd__o21ai_1
X_1698_ _2030_/A VGND VGND VPWR VPWR _1763_/A sky130_fd_sc_hd__clkbuf_2
X_3368_ _2520_/Y _2518_/Y _3374_/S VGND VGND VPWR VPWR _3368_/X sky130_fd_sc_hd__mux2_2
XFILLER_57_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2319_ _2263_/A _3096_/B _2294_/X _2640_/B VGND VGND VPWR VPWR _2319_/X sky130_fd_sc_hd__o22a_1
X_3299_ _1955_/Y _1950_/Y _3365_/S VGND VGND VPWR VPWR _3299_/X sky130_fd_sc_hd__mux2_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput21 _3156_/X VGND VGND VPWR VPWR output_thermometer_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput43 _3169_/X VGND VGND VPWR VPWR output_thermometer_o[41] sky130_fd_sc_hd__clkbuf_2
Xoutput32 _3271_/X VGND VGND VPWR VPWR output_thermometer_o[143] sky130_fd_sc_hd__clkbuf_2
Xoutput54 _3345_/X VGND VGND VPWR VPWR output_thermometer_o[217] sky130_fd_sc_hd__clkbuf_2
Xoutput65 _3207_/X VGND VGND VPWR VPWR output_thermometer_o[79] sky130_fd_sc_hd__clkbuf_2
Xoutput76 _3154_/X VGND VGND VPWR VPWR output_thermometer_o[26] sky130_fd_sc_hd__clkbuf_2
Xoutput87 _3180_/X VGND VGND VPWR VPWR output_thermometer_o[52] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput98 _3356_/X VGND VGND VPWR VPWR output_thermometer_o[228] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ _3126_/B _2611_/X _2406_/A _2097_/X VGND VGND VPWR VPWR _2670_/X sky130_fd_sc_hd__o22a_1
X_1621_ _2817_/A VGND VGND VPWR VPWR _2832_/A sky130_fd_sc_hd__buf_2
X_3222_ _2930_/Y _2928_/Y _3380_/S VGND VGND VPWR VPWR _3222_/X sky130_fd_sc_hd__mux2_1
X_3153_ _2678_/Y _2676_/Y _3346_/S VGND VGND VPWR VPWR _3153_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2104_ _3057_/A VGND VGND VPWR VPWR _2879_/C sky130_fd_sc_hd__buf_2
X_3084_ _3099_/A _3084_/B _3094_/C VGND VGND VPWR VPWR _3084_/X sky130_fd_sc_hd__or3_2
X_2035_ _2207_/A VGND VGND VPWR VPWR _2036_/A sky130_fd_sc_hd__inv_2
X_2937_ _2857_/X _1816_/B _2921_/X _2703_/B _2936_/X VGND VGND VPWR VPWR _2937_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2868_ _2886_/A _2868_/B VGND VGND VPWR VPWR _2868_/Y sky130_fd_sc_hd__nor2_1
X_2799_ _2920_/A VGND VGND VPWR VPWR _2799_/X sky130_fd_sc_hd__clkbuf_2
X_1819_ _1951_/A VGND VGND VPWR VPWR _1890_/A sky130_fd_sc_hd__buf_4
XFILLER_45_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2722_ _2737_/A _2722_/B VGND VGND VPWR VPWR _2722_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2653_ _2723_/A VGND VGND VPWR VPWR _2653_/X sky130_fd_sc_hd__buf_2
X_1604_ _1683_/A VGND VGND VPWR VPWR _1605_/B sky130_fd_sc_hd__buf_1
X_2584_ _2792_/B VGND VGND VPWR VPWR _2584_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3205_ _2870_/Y _2868_/Y _3330_/S VGND VGND VPWR VPWR _3205_/X sky130_fd_sc_hd__mux2_2
X_3136_ _2619_/Y _2617_/X _3351_/S VGND VGND VPWR VPWR _3136_/X sky130_fd_sc_hd__mux2_2
XFILLER_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3067_ _3110_/A VGND VGND VPWR VPWR _3083_/A sky130_fd_sc_hd__clkbuf_2
X_2018_ _2018_/A VGND VGND VPWR VPWR _2141_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2705_ _2705_/A _2936_/B VGND VGND VPWR VPWR _2705_/X sky130_fd_sc_hd__or2_1
X_2636_ _2636_/A _2636_/B VGND VGND VPWR VPWR _2636_/Y sky130_fd_sc_hd__nor2_1
Xoutput200 _3257_/X VGND VGND VPWR VPWR output_thermometer_o[129] sky130_fd_sc_hd__clkbuf_2
Xoutput233 _3381_/X VGND VGND VPWR VPWR output_thermometer_o[253] sky130_fd_sc_hd__clkbuf_2
Xoutput211 _3305_/X VGND VGND VPWR VPWR output_thermometer_o[177] sky130_fd_sc_hd__clkbuf_2
Xoutput244 _3254_/X VGND VGND VPWR VPWR output_thermometer_o[126] sky130_fd_sc_hd__clkbuf_2
Xoutput222 _3168_/X VGND VGND VPWR VPWR output_thermometer_o[40] sky130_fd_sc_hd__clkbuf_2
X_2567_ _1653_/X _3038_/B _2566_/X VGND VGND VPWR VPWR _2567_/Y sky130_fd_sc_hd__o21ai_1
Xoutput255 _3194_/X VGND VGND VPWR VPWR output_thermometer_o[66] sky130_fd_sc_hd__clkbuf_2
Xoutput266 _3355_/X VGND VGND VPWR VPWR output_thermometer_o[227] sky130_fd_sc_hd__clkbuf_2
X_2498_ _2741_/B _2483_/X _2497_/X VGND VGND VPWR VPWR _2498_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3119_ _3097_/X _2891_/B _3098_/X _2659_/B _3118_/X VGND VGND VPWR VPWR _3119_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2421_ _2421_/A VGND VGND VPWR VPWR _2421_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2352_ _1639_/X _2022_/A _2391_/A VGND VGND VPWR VPWR _2355_/A sky130_fd_sc_hd__o21ai_2
X_2283_ _2290_/A _3084_/B VGND VGND VPWR VPWR _2283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1998_ _2026_/A _1998_/B VGND VGND VPWR VPWR _2756_/B sky130_fd_sc_hd__nor2_2
X_2619_ _3074_/B _2602_/X _1610_/X _2271_/Y _2618_/X VGND VGND VPWR VPWR _2619_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2970_ _2970_/A VGND VGND VPWR VPWR _2985_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1921_ _1981_/A _2279_/A VGND VGND VPWR VPWR _1922_/A sky130_fd_sc_hd__or2_2
X_1852_ _1878_/A _1852_/B VGND VGND VPWR VPWR _1852_/Y sky130_fd_sc_hd__nor2_1
X_1783_ _1783_/A _3004_/A VGND VGND VPWR VPWR _1783_/X sky130_fd_sc_hd__or2_1
X_2404_ _2381_/X _2897_/B _2188_/X _3123_/B VGND VGND VPWR VPWR _2404_/X sky130_fd_sc_hd__o22a_1
X_3384_ _3408_/CLK input5/X VGND VGND VPWR VPWR _3384_/Q sky130_fd_sc_hd__dfxtp_2
X_2335_ _2335_/A VGND VGND VPWR VPWR _2335_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2266_ _2266_/A VGND VGND VPWR VPWR _2618_/A sky130_fd_sc_hd__inv_2
X_2197_ _2131_/X _2823_/B _2196_/X VGND VGND VPWR VPWR _2197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _3264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2120_ _2122_/B VGND VGND VPWR VPWR _3029_/B sky130_fd_sc_hd__inv_2
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2051_ _2081_/A _2051_/B VGND VGND VPWR VPWR _2772_/B sky130_fd_sc_hd__nor2_2
XFILLER_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2953_ _2956_/A _2953_/B VGND VGND VPWR VPWR _2953_/X sky130_fd_sc_hd__or2_1
X_1904_ _2082_/C VGND VGND VPWR VPWR _1954_/C sky130_fd_sc_hd__buf_1
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2884_ _2887_/A _3111_/B _3049_/C VGND VGND VPWR VPWR _2884_/X sky130_fd_sc_hd__or3_2
X_1835_ _1835_/A VGND VGND VPWR VPWR _2452_/A sky130_fd_sc_hd__inv_2
X_1766_ _2232_/A _1766_/B VGND VGND VPWR VPWR _2694_/B sky130_fd_sc_hd__nor2_2
X_1697_ _1581_/X _2676_/B _1696_/X VGND VGND VPWR VPWR _1697_/Y sky130_fd_sc_hd__o21ai_1
X_3367_ _2517_/Y _2515_/Y _3370_/S VGND VGND VPWR VPWR _3367_/X sky130_fd_sc_hd__mux2_4
X_2318_ _2318_/A _2344_/A VGND VGND VPWR VPWR _2640_/B sky130_fd_sc_hd__nor2_2
X_3298_ _1942_/Y _1938_/Y _3383_/S VGND VGND VPWR VPWR _3298_/X sky130_fd_sc_hd__mux2_2
X_2249_ _2249_/A VGND VGND VPWR VPWR _3068_/B sky130_fd_sc_hd__inv_2
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput22 _3147_/X VGND VGND VPWR VPWR output_thermometer_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput33 _3321_/X VGND VGND VPWR VPWR output_thermometer_o[193] sky130_fd_sc_hd__clkbuf_2
Xoutput66 _3272_/X VGND VGND VPWR VPWR output_thermometer_o[144] sky130_fd_sc_hd__clkbuf_2
Xoutput55 _3240_/X VGND VGND VPWR VPWR output_thermometer_o[112] sky130_fd_sc_hd__clkbuf_2
Xoutput44 _3131_/X VGND VGND VPWR VPWR output_thermometer_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput77 _3174_/X VGND VGND VPWR VPWR output_thermometer_o[46] sky130_fd_sc_hd__clkbuf_2
Xoutput99 _3358_/X VGND VGND VPWR VPWR output_thermometer_o[230] sky130_fd_sc_hd__clkbuf_2
Xoutput88 _3351_/X VGND VGND VPWR VPWR output_thermometer_o[223] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1620_ _2168_/B _2762_/A VGND VGND VPWR VPWR _2817_/A sky130_fd_sc_hd__or2_1
X_3221_ _2926_/Y _2924_/Y _3347_/S VGND VGND VPWR VPWR _3221_/X sky130_fd_sc_hd__mux2_2
X_3152_ _2675_/Y _2672_/Y _3382_/S VGND VGND VPWR VPWR _3152_/X sky130_fd_sc_hd__mux2_1
X_2103_ _2103_/A _2514_/B VGND VGND VPWR VPWR _2993_/B sky130_fd_sc_hd__or2_2
X_3083_ _3083_/A _3083_/B VGND VGND VPWR VPWR _3083_/Y sky130_fd_sc_hd__nor2_1
X_2034_ _2087_/A VGND VGND VPWR VPWR _2034_/X sky130_fd_sc_hd__buf_2
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2936_ _2936_/A _2936_/B VGND VGND VPWR VPWR _2936_/X sky130_fd_sc_hd__or2_1
X_2867_ _2867_/A VGND VGND VPWR VPWR _2886_/A sky130_fd_sc_hd__clkbuf_2
X_1818_ _1818_/A VGND VGND VPWR VPWR _1818_/X sky130_fd_sc_hd__buf_2
X_2798_ _2811_/A _2798_/B VGND VGND VPWR VPWR _2798_/Y sky130_fd_sc_hd__nor2_1
X_1749_ _1786_/A _2925_/A VGND VGND VPWR VPWR _1749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2721_ _2759_/A VGND VGND VPWR VPWR _2737_/A sky130_fd_sc_hd__clkbuf_2
X_2652_ _2659_/A _2652_/B VGND VGND VPWR VPWR _2652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1603_ _1624_/B _1791_/B VGND VGND VPWR VPWR _1683_/A sky130_fd_sc_hd__or2_4
X_2583_ _2589_/A VGND VGND VPWR VPWR _2792_/B sky130_fd_sc_hd__clkbuf_2
X_3204_ _2866_/Y _2864_/Y _3351_/S VGND VGND VPWR VPWR _3204_/X sky130_fd_sc_hd__mux2_2
X_3135_ _2616_/Y _2614_/X _3351_/S VGND VGND VPWR VPWR _3135_/X sky130_fd_sc_hd__mux2_2
X_3066_ _3052_/X _2839_/B _3053_/X _2605_/B _3065_/X VGND VGND VPWR VPWR _3066_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2017_ _2056_/A _2998_/B VGND VGND VPWR VPWR _2017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2919_ _2924_/A _2919_/B VGND VGND VPWR VPWR _2919_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2704_ _2723_/A VGND VGND VPWR VPWR _2704_/X sky130_fd_sc_hd__clkbuf_2
Xoutput201 _3198_/X VGND VGND VPWR VPWR output_thermometer_o[70] sky130_fd_sc_hd__clkbuf_2
X_2635_ _2606_/X _2864_/B _2634_/X VGND VGND VPWR VPWR _2635_/Y sky130_fd_sc_hd__o21ai_1
Xoutput234 _3199_/X VGND VGND VPWR VPWR output_thermometer_o[71] sky130_fd_sc_hd__clkbuf_2
Xoutput223 _3185_/X VGND VGND VPWR VPWR output_thermometer_o[57] sky130_fd_sc_hd__clkbuf_2
Xoutput212 _3359_/X VGND VGND VPWR VPWR output_thermometer_o[231] sky130_fd_sc_hd__clkbuf_2
Xoutput267 _3197_/X VGND VGND VPWR VPWR output_thermometer_o[69] sky130_fd_sc_hd__clkbuf_2
X_2566_ _2808_/B _2390_/X _3039_/B _2206_/X VGND VGND VPWR VPWR _2566_/X sky130_fd_sc_hd__o22a_1
Xoutput245 _3313_/X VGND VGND VPWR VPWR output_thermometer_o[185] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_clk_i clkbuf_0_clk_i/X VGND VGND VPWR VPWR _3404_/CLK sky130_fd_sc_hd__clkbuf_1
Xoutput256 _3286_/X VGND VGND VPWR VPWR output_thermometer_o[158] sky130_fd_sc_hd__clkbuf_2
X_2497_ _2478_/X _2974_/B _1950_/B _2488_/X VGND VGND VPWR VPWR _2497_/X sky130_fd_sc_hd__o22a_1
X_3118_ _3124_/A _3118_/B VGND VGND VPWR VPWR _3118_/X sky130_fd_sc_hd__or2_1
XFILLER_67_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3049_ _3058_/A _3049_/B _3049_/C VGND VGND VPWR VPWR _3049_/X sky130_fd_sc_hd__or3_2
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2420_ _2681_/B _2171_/X _2419_/X VGND VGND VPWR VPWR _2420_/Y sky130_fd_sc_hd__o21ai_1
X_2351_ _2682_/A VGND VGND VPWR VPWR _2351_/X sky130_fd_sc_hd__clkbuf_2
X_2282_ _2286_/A _2289_/B VGND VGND VPWR VPWR _3084_/B sky130_fd_sc_hd__nor2_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1997_ _1991_/A _1890_/A _1961_/X VGND VGND VPWR VPWR _2989_/B sky130_fd_sc_hd__a21oi_4
X_2618_ _2618_/A _2618_/B VGND VGND VPWR VPWR _2618_/X sky130_fd_sc_hd__or2_1
X_2549_ _2549_/A VGND VGND VPWR VPWR _2549_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1920_ _1920_/A VGND VGND VPWR VPWR _2279_/A sky130_fd_sc_hd__clkbuf_4
X_1851_ _1857_/B VGND VGND VPWR VPWR _1852_/B sky130_fd_sc_hd__inv_2
X_1782_ _2168_/A _2578_/A VGND VGND VPWR VPWR _3004_/A sky130_fd_sc_hd__or2_4
X_2403_ _2403_/A VGND VGND VPWR VPWR _3123_/B sky130_fd_sc_hd__inv_2
X_3383_ _2573_/X _3383_/A1 _3383_/S VGND VGND VPWR VPWR _3383_/X sky130_fd_sc_hd__mux2_1
X_2334_ _2334_/A VGND VGND VPWR VPWR _2335_/A sky130_fd_sc_hd__buf_1
X_2265_ _2265_/A _2265_/B _2268_/B VGND VGND VPWR VPWR _2266_/A sky130_fd_sc_hd__or3_4
X_2196_ _2188_/X _3048_/B _2606_/A _2588_/B VGND VGND VPWR VPWR _2196_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 _3338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2050_ _1992_/X _2019_/X _2020_/X _2530_/A _2023_/X VGND VGND VPWR VPWR _3003_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_19_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2952_ _2967_/A _2952_/B VGND VGND VPWR VPWR _2952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1903_ _1903_/A _1903_/B VGND VGND VPWR VPWR _2726_/B sky130_fd_sc_hd__nor2_4
X_2883_ _3057_/A VGND VGND VPWR VPWR _3049_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1834_ _2067_/A _2029_/A VGND VGND VPWR VPWR _1835_/A sky130_fd_sc_hd__or2_2
X_1765_ _1786_/A _2929_/A VGND VGND VPWR VPWR _1765_/Y sky130_fd_sc_hd__nor2_1
X_1696_ _1610_/X _2413_/A _1622_/X _2910_/B VGND VGND VPWR VPWR _1696_/X sky130_fd_sc_hd__o22a_1
X_3366_ _2513_/Y _2510_/Y _3370_/S VGND VGND VPWR VPWR _3366_/X sky130_fd_sc_hd__mux2_2
X_3297_ _1930_/Y _1925_/Y _3365_/S VGND VGND VPWR VPWR _3297_/X sky130_fd_sc_hd__mux2_2
X_2317_ _2318_/A _2317_/B VGND VGND VPWR VPWR _3096_/B sky130_fd_sc_hd__nor2_2
X_2248_ _2549_/A VGND VGND VPWR VPWR _2248_/X sky130_fd_sc_hd__clkbuf_2
X_2179_ _2189_/B VGND VGND VPWR VPWR _2338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput34 _3357_/X VGND VGND VPWR VPWR output_thermometer_o[229] sky130_fd_sc_hd__clkbuf_2
Xoutput23 _3256_/X VGND VGND VPWR VPWR output_thermometer_o[128] sky130_fd_sc_hd__clkbuf_2
Xoutput56 _3284_/X VGND VGND VPWR VPWR output_thermometer_o[156] sky130_fd_sc_hd__clkbuf_2
Xoutput67 _3278_/X VGND VGND VPWR VPWR output_thermometer_o[150] sky130_fd_sc_hd__clkbuf_2
Xoutput45 _3167_/X VGND VGND VPWR VPWR output_thermometer_o[39] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput89 _3153_/X VGND VGND VPWR VPWR output_thermometer_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput78 _3139_/X VGND VGND VPWR VPWR output_thermometer_o[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3220_ _2923_/Y _2919_/Y _3380_/S VGND VGND VPWR VPWR _3220_/X sky130_fd_sc_hd__mux2_1
X_3151_ _2671_/Y _2669_/Y _3382_/S VGND VGND VPWR VPWR _3151_/X sky130_fd_sc_hd__mux2_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2102_ _2265_/B _1570_/A _2101_/Y VGND VGND VPWR VPWR _2514_/B sky130_fd_sc_hd__o21ai_2
X_3082_ _3078_/X _2853_/B _3079_/X _2621_/B _3081_/X VGND VGND VPWR VPWR _3082_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2033_ _2056_/A _3001_/B VGND VGND VPWR VPWR _2033_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ _2948_/A _2935_/B VGND VGND VPWR VPWR _2935_/Y sky130_fd_sc_hd__nor2_1
X_2866_ _1818_/X _2633_/B _2865_/X VGND VGND VPWR VPWR _2866_/Y sky130_fd_sc_hd__o21ai_1
X_1817_ _2817_/A VGND VGND VPWR VPWR _1818_/A sky130_fd_sc_hd__clkbuf_2
X_2797_ _2867_/A VGND VGND VPWR VPWR _2811_/A sky130_fd_sc_hd__clkbuf_2
X_1748_ _1752_/B VGND VGND VPWR VPWR _2925_/A sky130_fd_sc_hd__inv_2
X_1679_ _1566_/A _1847_/A _1584_/A VGND VGND VPWR VPWR _1808_/B sky130_fd_sc_hd__o21ai_4
X_3349_ _2433_/Y _2431_/Y _3380_/S VGND VGND VPWR VPWR _3349_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2720_ _1878_/B _2704_/X _2952_/B _2715_/X _2719_/X VGND VGND VPWR VPWR _2720_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2651_ _3107_/B _2630_/X _2626_/X _2878_/B _2650_/X VGND VGND VPWR VPWR _2651_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1602_ _2178_/A _1860_/A _1570_/A _3390_/Q VGND VGND VPWR VPWR _1791_/B sky130_fd_sc_hd__o31a_1
X_2582_ _2815_/A _2582_/B VGND VGND VPWR VPWR _2589_/A sky130_fd_sc_hd__or2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3203_ _2863_/Y _2861_/Y _3330_/S VGND VGND VPWR VPWR _3203_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3134_ _2613_/Y _2610_/Y _3342_/S VGND VGND VPWR VPWR _3134_/X sky130_fd_sc_hd__mux2_2
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3065_ _3108_/A _3065_/B VGND VGND VPWR VPWR _3065_/X sky130_fd_sc_hd__or2_1
XFILLER_67_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2016_ _2026_/B VGND VGND VPWR VPWR _2998_/B sky130_fd_sc_hd__inv_2
X_2918_ _1725_/C _2901_/X _2872_/X _2685_/B _2917_/X VGND VGND VPWR VPWR _2918_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2849_ _2849_/A VGND VGND VPWR VPWR _2849_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2703_ _2718_/A _2703_/B VGND VGND VPWR VPWR _2703_/Y sky130_fd_sc_hd__nor2_1
X_2634_ _2341_/X _3090_/A _2299_/B _2584_/X VGND VGND VPWR VPWR _2634_/X sky130_fd_sc_hd__o22a_1
Xoutput235 _3309_/X VGND VGND VPWR VPWR output_thermometer_o[181] sky130_fd_sc_hd__clkbuf_2
X_2565_ _2565_/A _2809_/A VGND VGND VPWR VPWR _2565_/Y sky130_fd_sc_hd__nor2_1
Xoutput213 _3173_/X VGND VGND VPWR VPWR output_thermometer_o[45] sky130_fd_sc_hd__clkbuf_2
Xoutput224 _3136_/X VGND VGND VPWR VPWR output_thermometer_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput202 _3166_/X VGND VGND VPWR VPWR output_thermometer_o[38] sky130_fd_sc_hd__clkbuf_2
Xoutput246 _3369_/X VGND VGND VPWR VPWR output_thermometer_o[241] sky130_fd_sc_hd__clkbuf_2
Xoutput257 _3326_/X VGND VGND VPWR VPWR output_thermometer_o[198] sky130_fd_sc_hd__clkbuf_2
Xoutput268 _3383_/X VGND VGND VPWR VPWR output_thermometer_o[255] sky130_fd_sc_hd__clkbuf_2
X_2496_ _2975_/B VGND VGND VPWR VPWR _2496_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3117_ _3126_/A _3117_/B VGND VGND VPWR VPWR _3117_/Y sky130_fd_sc_hd__nor2_1
X_3048_ _3064_/A _3048_/B VGND VGND VPWR VPWR _3048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2350_ _3108_/B VGND VGND VPWR VPWR _2350_/Y sky130_fd_sc_hd__inv_2
X_2281_ _2212_/X _2853_/B _2280_/X VGND VGND VPWR VPWR _2281_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ _1996_/A _1996_/B VGND VGND VPWR VPWR _1996_/Y sky130_fd_sc_hd__nor2_1
X_2617_ _2617_/A _2617_/B VGND VGND VPWR VPWR _2617_/X sky130_fd_sc_hd__or2_1
X_2548_ _2548_/A _2548_/B VGND VGND VPWR VPWR _2548_/Y sky130_fd_sc_hd__nor2_1
X_2479_ _2478_/X _2958_/B _1899_/B _2464_/X VGND VGND VPWR VPWR _2479_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1850_ _1806_/X _2457_/A _2093_/A VGND VGND VPWR VPWR _1857_/B sky130_fd_sc_hd__o21ai_2
X_1781_ _2837_/A _1783_/A VGND VGND VPWR VPWR _2931_/B sky130_fd_sc_hd__and2_1
X_3382_ _2570_/Y _2568_/Y _3382_/S VGND VGND VPWR VPWR _3382_/X sky130_fd_sc_hd__mux2_2
X_2402_ _2184_/A _2398_/B _2142_/A VGND VGND VPWR VPWR _2897_/B sky130_fd_sc_hd__o21a_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2333_ _2333_/A _2333_/B VGND VGND VPWR VPWR _2334_/A sky130_fd_sc_hd__or2_1
X_2264_ _2256_/X _2258_/Y _2080_/X _2848_/B _2263_/X VGND VGND VPWR VPWR _2264_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2195_ _2195_/A _2286_/B VGND VGND VPWR VPWR _2588_/B sky130_fd_sc_hd__nor2_2
XFILLER_25_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1979_ _1974_/X _2982_/B _1963_/X _2749_/B _1978_/X VGND VGND VPWR VPWR _1979_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 _3215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2951_ _2970_/A VGND VGND VPWR VPWR _2967_/A sky130_fd_sc_hd__clkbuf_2
X_1902_ _2025_/A VGND VGND VPWR VPWR _1902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2882_ _3097_/A VGND VGND VPWR VPWR _2882_/X sky130_fd_sc_hd__buf_2
X_1833_ _1833_/A _2057_/A VGND VGND VPWR VPWR _2029_/A sky130_fd_sc_hd__or2_1
X_1764_ _1766_/B VGND VGND VPWR VPWR _2929_/A sky130_fd_sc_hd__inv_2
X_1695_ _1725_/A _1725_/B _1695_/C VGND VGND VPWR VPWR _2910_/B sky130_fd_sc_hd__and3_1
X_3365_ _2508_/Y _2505_/Y _3365_/S VGND VGND VPWR VPWR _3365_/X sky130_fd_sc_hd__mux2_4
X_2316_ _2291_/X _3099_/B _2837_/A VGND VGND VPWR VPWR _2871_/B sky130_fd_sc_hd__o21a_1
XFILLER_57_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3296_ _1918_/Y _1912_/Y _3383_/S VGND VGND VPWR VPWR _3296_/X sky130_fd_sc_hd__mux2_1
X_2247_ _2233_/X _2240_/B _2234_/X VGND VGND VPWR VPWR _2845_/B sky130_fd_sc_hd__o21a_1
X_2178_ _2178_/A _2178_/B VGND VGND VPWR VPWR _2189_/B sky130_fd_sc_hd__or2_2
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput24 _3273_/X VGND VGND VPWR VPWR output_thermometer_o[145] sky130_fd_sc_hd__clkbuf_2
Xoutput13 _3392_/Q VGND VGND VPWR VPWR output_binary_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput46 _3146_/X VGND VGND VPWR VPWR output_thermometer_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput57 _3317_/X VGND VGND VPWR VPWR output_thermometer_o[189] sky130_fd_sc_hd__clkbuf_2
Xoutput35 _3195_/X VGND VGND VPWR VPWR output_thermometer_o[67] sky130_fd_sc_hd__clkbuf_2
Xoutput79 _3216_/X VGND VGND VPWR VPWR output_thermometer_o[88] sky130_fd_sc_hd__clkbuf_2
Xoutput68 _3265_/X VGND VGND VPWR VPWR output_thermometer_o[137] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3150_ _2668_/Y _2666_/Y _3342_/S VGND VGND VPWR VPWR _3150_/X sky130_fd_sc_hd__mux2_2
X_2101_ _2101_/A _2161_/A VGND VGND VPWR VPWR _2101_/Y sky130_fd_sc_hd__nor2_2
XFILLER_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3081_ _3099_/A _3081_/B _3094_/C VGND VGND VPWR VPWR _3081_/X sky130_fd_sc_hd__or3_2
X_2032_ _2039_/B VGND VGND VPWR VPWR _3001_/B sky130_fd_sc_hd__inv_2
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2934_ _1858_/A _2854_/B _2301_/A _2821_/B _2173_/X VGND VGND VPWR VPWR _2934_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2865_ _3054_/A _3090_/A _2331_/X _3091_/B VGND VGND VPWR VPWR _2865_/X sky130_fd_sc_hd__o22a_1
X_1816_ _1878_/A _1816_/B VGND VGND VPWR VPWR _1816_/Y sky130_fd_sc_hd__nor2_1
X_2796_ _3025_/B _2761_/X _3024_/B _2791_/X _2795_/X VGND VGND VPWR VPWR _2796_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1747_ _1763_/A _1747_/B _1747_/C VGND VGND VPWR VPWR _1752_/B sky130_fd_sc_hd__or3_4
X_1678_ _3384_/Q VGND VGND VPWR VPWR _1809_/B sky130_fd_sc_hd__inv_2
X_3348_ _2430_/Y _2425_/Y _3380_/S VGND VGND VPWR VPWR _3348_/X sky130_fd_sc_hd__mux2_2
X_3279_ _1634_/Y _3126_/Y _3342_/S VGND VGND VPWR VPWR _3279_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2650_ _2650_/A _2660_/B VGND VGND VPWR VPWR _2650_/X sky130_fd_sc_hd__or2_1
X_1601_ _1601_/A VGND VGND VPWR VPWR _1624_/B sky130_fd_sc_hd__inv_2
X_2581_ _2581_/A VGND VGND VPWR VPWR _2581_/X sky130_fd_sc_hd__clkbuf_2
X_3202_ _2860_/Y _2856_/Y _3330_/S VGND VGND VPWR VPWR _3202_/X sky130_fd_sc_hd__mux2_2
X_3133_ _2609_/Y _2605_/Y _3342_/S VGND VGND VPWR VPWR _3133_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3064_ _3064_/A _3064_/B VGND VGND VPWR VPWR _3064_/Y sky130_fd_sc_hd__nor2_1
X_2015_ _2005_/X _2195_/A _2397_/A _2014_/X VGND VGND VPWR VPWR _2026_/B sky130_fd_sc_hd__a31o_1
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2917_ _2917_/A _2922_/B VGND VGND VPWR VPWR _2917_/X sky130_fd_sc_hd__or2_1
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2848_ _2931_/A _2848_/B VGND VGND VPWR VPWR _2848_/Y sky130_fd_sc_hd__nor2_1
X_2779_ _2889_/A VGND VGND VPWR VPWR _2867_/A sky130_fd_sc_hd__buf_2
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2702_ _2759_/A VGND VGND VPWR VPWR _2718_/A sky130_fd_sc_hd__clkbuf_2
X_2633_ _2636_/A _2633_/B VGND VGND VPWR VPWR _2633_/Y sky130_fd_sc_hd__nor2_1
Xoutput214 _3382_/X VGND VGND VPWR VPWR output_thermometer_o[254] sky130_fd_sc_hd__clkbuf_2
Xoutput225 _3178_/X VGND VGND VPWR VPWR output_thermometer_o[50] sky130_fd_sc_hd__clkbuf_2
Xoutput203 _3315_/X VGND VGND VPWR VPWR output_thermometer_o[187] sky130_fd_sc_hd__clkbuf_2
X_2564_ _2805_/B _2545_/X _2563_/X VGND VGND VPWR VPWR _2564_/Y sky130_fd_sc_hd__o21ai_1
Xoutput247 _3348_/X VGND VGND VPWR VPWR output_thermometer_o[220] sky130_fd_sc_hd__clkbuf_2
Xoutput236 _3235_/X VGND VGND VPWR VPWR output_thermometer_o[107] sky130_fd_sc_hd__clkbuf_2
Xoutput258 _3159_/X VGND VGND VPWR VPWR output_thermometer_o[31] sky130_fd_sc_hd__clkbuf_2
Xoutput269 _3342_/X VGND VGND VPWR VPWR output_thermometer_o[214] sky130_fd_sc_hd__clkbuf_2
X_2495_ _2495_/A _2495_/B VGND VGND VPWR VPWR _2975_/B sky130_fd_sc_hd__or2_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3116_ _3097_/X _2886_/B _3098_/X _2656_/B _3115_/X VGND VGND VPWR VPWR _3116_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_55_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3047_ _3047_/A VGND VGND VPWR VPWR _3064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2280_ _2188_/X _3077_/B _2606_/A _2621_/B VGND VGND VPWR VPWR _2280_/X sky130_fd_sc_hd__o22a_1
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1995_ _1998_/B VGND VGND VPWR VPWR _1996_/B sky130_fd_sc_hd__inv_2
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2616_ _3071_/B _2602_/X _2594_/X _2848_/B _2615_/X VGND VGND VPWR VPWR _2616_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2547_ _2787_/B _2545_/X _2546_/X VGND VGND VPWR VPWR _2547_/Y sky130_fd_sc_hd__o21ai_1
X_2478_ _2478_/A VGND VGND VPWR VPWR _2478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1780_ _2932_/A _2018_/A VGND VGND VPWR VPWR _1783_/A sky130_fd_sc_hd__or2_1
X_3381_ _2567_/Y _2565_/Y _3381_/S VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__mux2_1
X_2401_ _2401_/A _2403_/A VGND VGND VPWR VPWR _2666_/B sky130_fd_sc_hd__nor2_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2332_ _2265_/A _2265_/B _2165_/B VGND VGND VPWR VPWR _2333_/B sky130_fd_sc_hd__o21a_1
X_2263_ _2263_/A _3071_/B VGND VGND VPWR VPWR _2263_/X sky130_fd_sc_hd__or2_1
X_2194_ _2344_/A VGND VGND VPWR VPWR _2286_/B sky130_fd_sc_hd__buf_2
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1978_ _1978_/A _2504_/A _2071_/C VGND VGND VPWR VPWR _1978_/X sky130_fd_sc_hd__or3_1
XFILLER_68_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2950_ _2940_/X _1865_/B _2941_/X _2714_/B _2949_/X VGND VGND VPWR VPWR _2950_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2881_ _2886_/A _2881_/B VGND VGND VPWR VPWR _2881_/Y sky130_fd_sc_hd__nor2_1
X_1901_ _1890_/X _2252_/B _1900_/X VGND VGND VPWR VPWR _2958_/B sky130_fd_sc_hd__a21oi_4
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1832_ _1832_/A VGND VGND VPWR VPWR _2057_/A sky130_fd_sc_hd__clkbuf_2
X_1763_ _1763_/A _1763_/B _2044_/A VGND VGND VPWR VPWR _1766_/B sky130_fd_sc_hd__or3_4
X_1694_ _1769_/A _1695_/C VGND VGND VPWR VPWR _2413_/A sky130_fd_sc_hd__or2_2
X_3364_ _2503_/Y _2500_/Y _3365_/S VGND VGND VPWR VPWR _3364_/X sky130_fd_sc_hd__mux2_2
X_2315_ _2315_/A VGND VGND VPWR VPWR _2315_/X sky130_fd_sc_hd__buf_2
X_3295_ _1906_/Y _1899_/Y _3365_/S VGND VGND VPWR VPWR _3295_/X sky130_fd_sc_hd__mux2_2
XFILLER_57_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2246_ _2478_/A VGND VGND VPWR VPWR _2246_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2177_ _3058_/A VGND VGND VPWR VPWR _2290_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput25 _3171_/X VGND VGND VPWR VPWR output_thermometer_o[43] sky130_fd_sc_hd__clkbuf_2
Xoutput14 _3393_/Q VGND VGND VPWR VPWR output_binary_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput36 _3304_/X VGND VGND VPWR VPWR output_thermometer_o[176] sky130_fd_sc_hd__clkbuf_2
Xoutput47 _3205_/X VGND VGND VPWR VPWR output_thermometer_o[77] sky130_fd_sc_hd__clkbuf_2
Xoutput58 _3324_/X VGND VGND VPWR VPWR output_thermometer_o[196] sky130_fd_sc_hd__clkbuf_2
Xoutput69 _3211_/X VGND VGND VPWR VPWR output_thermometer_o[83] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2100_ _3027_/A _2100_/B VGND VGND VPWR VPWR _3021_/A sky130_fd_sc_hd__or2_2
X_3080_ _3080_/A VGND VGND VPWR VPWR _3099_/A sky130_fd_sc_hd__buf_1
X_2031_ _2005_/X _2207_/A _2030_/X _2014_/X VGND VGND VPWR VPWR _2039_/B sky130_fd_sc_hd__a31o_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2933_ _2440_/A _2825_/X _2921_/X _2697_/B _2932_/X VGND VGND VPWR VPWR _2933_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2864_ _2864_/A _2864_/B VGND VGND VPWR VPWR _2864_/Y sky130_fd_sc_hd__nor2_1
X_2795_ _2795_/A _2803_/B VGND VGND VPWR VPWR _2795_/X sky130_fd_sc_hd__or2_1
X_1815_ _1823_/B VGND VGND VPWR VPWR _1816_/B sky130_fd_sc_hd__inv_2
X_1746_ _2149_/B VGND VGND VPWR VPWR _1747_/B sky130_fd_sc_hd__inv_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1677_ _1691_/A VGND VGND VPWR VPWR _1684_/A sky130_fd_sc_hd__clkbuf_2
X_3347_ _2424_/Y _2421_/Y _3347_/S VGND VGND VPWR VPWR _3347_/X sky130_fd_sc_hd__mux2_1
X_3278_ _3125_/Y _3123_/Y _3342_/S VGND VGND VPWR VPWR _3278_/X sky130_fd_sc_hd__mux2_2
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2229_ _2359_/A _2229_/B VGND VGND VPWR VPWR _3065_/B sky130_fd_sc_hd__or2_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1600_ _2090_/A _2347_/A _2092_/C VGND VGND VPWR VPWR _1631_/A sky130_fd_sc_hd__o21ai_2
X_2580_ _2766_/A VGND VGND VPWR VPWR _2581_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3201_ _2855_/Y _2853_/Y _3330_/S VGND VGND VPWR VPWR _3201_/X sky130_fd_sc_hd__mux2_2
X_3132_ _2604_/Y _2600_/Y _3346_/S VGND VGND VPWR VPWR _3132_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3063_ _3052_/X _2836_/B _3053_/X _2600_/B _3062_/X VGND VGND VPWR VPWR _3063_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2014_ _2044_/A VGND VGND VPWR VPWR _2014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2916_ _2924_/A _2916_/B VGND VGND VPWR VPWR _2916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2847_ _2087_/X _2610_/B _2840_/X _3069_/B _2846_/X VGND VGND VPWR VPWR _2847_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2778_ _2534_/A _2763_/X _3008_/B _2773_/X _2777_/X VGND VGND VPWR VPWR _2778_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1729_ _1808_/B VGND VGND VPWR VPWR _1759_/A sky130_fd_sc_hd__inv_2
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2701_ _2301_/A _2581_/X _2700_/X VGND VGND VPWR VPWR _2701_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2632_ _3087_/B _2630_/X _2626_/X _2861_/B _2631_/X VGND VGND VPWR VPWR _2632_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput215 _3289_/X VGND VGND VPWR VPWR output_thermometer_o[161] sky130_fd_sc_hd__clkbuf_2
X_2563_ _1653_/A _3035_/B _3036_/B _2549_/X VGND VGND VPWR VPWR _2563_/X sky130_fd_sc_hd__o22a_1
Xoutput226 _3164_/X VGND VGND VPWR VPWR output_thermometer_o[36] sky130_fd_sc_hd__clkbuf_2
Xoutput204 _3151_/X VGND VGND VPWR VPWR output_thermometer_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput237 _3362_/X VGND VGND VPWR VPWR output_thermometer_o[234] sky130_fd_sc_hd__clkbuf_2
Xoutput259 _3312_/X VGND VGND VPWR VPWR output_thermometer_o[184] sky130_fd_sc_hd__clkbuf_2
Xoutput248 _3371_/X VGND VGND VPWR VPWR output_thermometer_o[243] sky130_fd_sc_hd__clkbuf_2
X_2494_ _2737_/B _2483_/X _2493_/X VGND VGND VPWR VPWR _2494_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3115_ _3124_/A _3115_/B VGND VGND VPWR VPWR _3115_/X sky130_fd_sc_hd__or2_1
X_3046_ _1789_/X _1792_/Y _1581_/X _3105_/A VGND VGND VPWR VPWR _3046_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ _2514_/A _1992_/X _2291_/A VGND VGND VPWR VPWR _1998_/B sky130_fd_sc_hd__o21ai_2
XFILLER_60_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2615_ _2705_/A _2615_/B VGND VGND VPWR VPWR _2615_/X sky130_fd_sc_hd__or2_1
X_2546_ _1653_/A _3018_/B _2086_/B _2531_/X VGND VGND VPWR VPWR _2546_/X sky130_fd_sc_hd__o22a_1
X_2477_ _2962_/B VGND VGND VPWR VPWR _2477_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3029_ _3029_/A _3029_/B VGND VGND VPWR VPWR _3029_/X sky130_fd_sc_hd__or2_1
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ _2400_/A _2400_/B VGND VGND VPWR VPWR _2403_/A sky130_fd_sc_hd__or2_2
X_3380_ _2564_/Y _2562_/Y _3380_/S VGND VGND VPWR VPWR _3380_/X sky130_fd_sc_hd__mux2_1
X_2331_ _2990_/A VGND VGND VPWR VPWR _2331_/X sky130_fd_sc_hd__buf_2
X_2262_ _2262_/A VGND VGND VPWR VPWR _3071_/B sky130_fd_sc_hd__inv_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2193_ _2193_/A _2277_/A VGND VGND VPWR VPWR _2344_/A sky130_fd_sc_hd__or2_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1977_ _2026_/A _1977_/B VGND VGND VPWR VPWR _2749_/B sky130_fd_sc_hd__nor2_2
X_2529_ _2769_/B _2527_/X _2528_/X VGND VGND VPWR VPWR _2529_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1900_ _1900_/A VGND VGND VPWR VPWR _1900_/X sky130_fd_sc_hd__buf_4
X_2880_ _2087_/X _2649_/B _2840_/X _3108_/B _2879_/X VGND VGND VPWR VPWR _2880_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1831_ _1818_/X _2935_/B _1777_/X _2703_/B _1830_/X VGND VGND VPWR VPWR _1831_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1762_ _2157_/B VGND VGND VPWR VPWR _1763_/B sky130_fd_sc_hd__inv_2
X_1693_ _2386_/A _1684_/B _1631_/B VGND VGND VPWR VPWR _1695_/C sky130_fd_sc_hd__o21ai_1
X_3363_ _2498_/Y _2496_/Y _3365_/S VGND VGND VPWR VPWR _3363_/X sky130_fd_sc_hd__mux2_1
X_2314_ _3058_/A _3099_/B VGND VGND VPWR VPWR _2314_/Y sky130_fd_sc_hd__nor2_1
X_3294_ _1894_/Y _1889_/Y _3383_/S VGND VGND VPWR VPWR _3294_/X sky130_fd_sc_hd__mux2_1
X_2245_ _2245_/A VGND VGND VPWR VPWR _2478_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2176_ _3080_/A VGND VGND VPWR VPWR _3058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput15 _3380_/X VGND VGND VPWR VPWR output_thermometer_o[252] sky130_fd_sc_hd__clkbuf_2
Xoutput26 _3367_/X VGND VGND VPWR VPWR output_thermometer_o[239] sky130_fd_sc_hd__clkbuf_2
Xoutput37 _3253_/X VGND VGND VPWR VPWR output_thermometer_o[125] sky130_fd_sc_hd__clkbuf_2
Xoutput48 _3377_/X VGND VGND VPWR VPWR output_thermometer_o[249] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput59 _3280_/X VGND VGND VPWR VPWR output_thermometer_o[152] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2030_ _2030_/A VGND VGND VPWR VPWR _2030_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2932_ _2932_/A _2932_/B VGND VGND VPWR VPWR _2932_/X sky130_fd_sc_hd__or2_1
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2863_ _2857_/X _3087_/B _2833_/X _2629_/B _2862_/X VGND VGND VPWR VPWR _2863_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2794_ _2794_/A _2794_/B VGND VGND VPWR VPWR _2794_/Y sky130_fd_sc_hd__nor2_1
X_1814_ _1806_/X _2446_/A _2093_/A VGND VGND VPWR VPWR _1823_/B sky130_fd_sc_hd__o21ai_2
X_1745_ _1761_/A _1968_/A VGND VGND VPWR VPWR _2149_/B sky130_fd_sc_hd__or2_4
X_1676_ _1653_/X _2672_/B _1660_/X _2905_/B _1675_/X VGND VGND VPWR VPWR _1676_/Y
+ sky130_fd_sc_hd__o221ai_2
X_3346_ _2420_/Y _2418_/Y _3346_/S VGND VGND VPWR VPWR _3346_/X sky130_fd_sc_hd__mux2_2
X_3277_ _3122_/Y _3120_/Y _3382_/S VGND VGND VPWR VPWR _3277_/X sky130_fd_sc_hd__mux2_1
X_2228_ _2239_/A _2231_/B VGND VGND VPWR VPWR _2229_/B sky130_fd_sc_hd__nor2_1
X_2159_ _1818_/A _3041_/B _2157_/B _1802_/A VGND VGND VPWR VPWR _2159_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3200_ _2852_/Y _2271_/A _3351_/S VGND VGND VPWR VPWR _3200_/X sky130_fd_sc_hd__mux2_2
X_3131_ _2599_/Y _2597_/Y _3346_/S VGND VGND VPWR VPWR _3131_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3062_ _3108_/A _3062_/B VGND VGND VPWR VPWR _3062_/X sky130_fd_sc_hd__or2_1
X_2013_ _2030_/A VGND VGND VPWR VPWR _2397_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2915_ _1712_/C _2901_/X _2872_/X _2681_/B _2914_/X VGND VGND VPWR VPWR _2915_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2846_ _2887_/A _3068_/B _2879_/C VGND VGND VPWR VPWR _2846_/X sky130_fd_sc_hd__or3_2
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2777_ _3009_/B _2782_/B VGND VGND VPWR VPWR _2777_/X sky130_fd_sc_hd__or2_1
X_1728_ _2568_/A VGND VGND VPWR VPWR _1786_/A sky130_fd_sc_hd__buf_2
X_1659_ _2832_/A VGND VGND VPWR VPWR _3097_/A sky130_fd_sc_hd__buf_1
XFILLER_58_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3329_ _2281_/Y _2275_/Y _3330_/S VGND VGND VPWR VPWR _3329_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2700_ _3054_/A _1794_/Y _1858_/A _2618_/B VGND VGND VPWR VPWR _2700_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2631_ _3088_/B _2641_/B VGND VGND VPWR VPWR _2631_/X sky130_fd_sc_hd__or2_1
X_2562_ _2565_/A _2806_/A VGND VGND VPWR VPWR _2562_/Y sky130_fd_sc_hd__nor2_1
Xoutput205 _3352_/X VGND VGND VPWR VPWR output_thermometer_o[224] sky130_fd_sc_hd__clkbuf_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput216 _3366_/X VGND VGND VPWR VPWR output_thermometer_o[238] sky130_fd_sc_hd__clkbuf_2
Xoutput227 _3338_/X VGND VGND VPWR VPWR output_thermometer_o[210] sky130_fd_sc_hd__clkbuf_2
Xoutput249 _3215_/X VGND VGND VPWR VPWR output_thermometer_o[87] sky130_fd_sc_hd__clkbuf_2
Xoutput238 _3145_/X VGND VGND VPWR VPWR output_thermometer_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2493_ _2478_/X _2971_/B _1938_/B _2488_/X VGND VGND VPWR VPWR _2493_/X sky130_fd_sc_hd__o22a_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3114_ _3126_/A _3114_/B VGND VGND VPWR VPWR _3114_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3045_ _3102_/A _2161_/Y _2577_/A _2166_/X VGND VGND VPWR VPWR _3045_/X sky130_fd_sc_hd__o211a_1
XFILLER_23_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2829_ _2936_/A _3054_/B VGND VGND VPWR VPWR _2829_/X sky130_fd_sc_hd__or2_1
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1993_ _2157_/C VGND VGND VPWR VPWR _2291_/A sky130_fd_sc_hd__buf_4
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2614_ _3387_/Q _2617_/B VGND VGND VPWR VPWR _2614_/X sky130_fd_sc_hd__or2_1
X_2545_ _2682_/A VGND VGND VPWR VPWR _2545_/X sky130_fd_sc_hd__buf_2
X_2476_ _2476_/A _2495_/B VGND VGND VPWR VPWR _2962_/B sky130_fd_sc_hd__or2_2
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3028_ _3041_/A _3028_/B VGND VGND VPWR VPWR _3028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2330_ _2993_/A VGND VGND VPWR VPWR _2990_/A sky130_fd_sc_hd__clkbuf_2
X_2261_ _2435_/A VGND VGND VPWR VPWR _2263_/A sky130_fd_sc_hd__buf_2
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2192_ _2390_/A VGND VGND VPWR VPWR _2606_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1976_ _2038_/A VGND VGND VPWR VPWR _2026_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2528_ _2523_/X _3000_/B _3001_/B _2511_/X VGND VGND VPWR VPWR _2528_/X sky130_fd_sc_hd__o22a_1
X_2459_ _2527_/A VGND VGND VPWR VPWR _2459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1830_ _1858_/A _2446_/A _3105_/A VGND VGND VPWR VPWR _1830_/X sky130_fd_sc_hd__or3_2
X_1761_ _1761_/A _1980_/A VGND VGND VPWR VPWR _2157_/B sky130_fd_sc_hd__or2_4
XFILLER_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1692_ _2030_/A VGND VGND VPWR VPWR _2386_/A sky130_fd_sc_hd__clkbuf_2
X_3362_ _2494_/Y _2492_/Y _3365_/S VGND VGND VPWR VPWR _3362_/X sky130_fd_sc_hd__mux2_2
X_2313_ _2318_/A _2338_/A VGND VGND VPWR VPWR _3099_/B sky130_fd_sc_hd__nor2_2
X_3293_ _1882_/Y _1878_/Y _3357_/S VGND VGND VPWR VPWR _3293_/X sky130_fd_sc_hd__mux2_1
X_2244_ _2380_/A _2249_/A VGND VGND VPWR VPWR _2610_/B sky130_fd_sc_hd__nor2_4
X_2175_ _2815_/A VGND VGND VPWR VPWR _3080_/A sky130_fd_sc_hd__buf_2
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1959_ _1964_/B VGND VGND VPWR VPWR _1960_/B sky130_fd_sc_hd__inv_2
Xoutput38 _3187_/X VGND VGND VPWR VPWR output_thermometer_o[59] sky130_fd_sc_hd__clkbuf_2
Xoutput27 _3196_/X VGND VGND VPWR VPWR output_thermometer_o[68] sky130_fd_sc_hd__clkbuf_2
Xoutput49 _3162_/X VGND VGND VPWR VPWR output_thermometer_o[34] sky130_fd_sc_hd__clkbuf_2
Xoutput16 _3157_/X VGND VGND VPWR VPWR output_thermometer_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2931_ _2931_/A _2931_/B VGND VGND VPWR VPWR _2931_/Y sky130_fd_sc_hd__nor2_1
X_2862_ _3088_/B _2932_/B VGND VGND VPWR VPWR _2862_/X sky130_fd_sc_hd__or2_1
X_2793_ _2095_/B _2761_/X _2100_/B _2791_/X _2792_/X VGND VGND VPWR VPWR _2793_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1813_ _2233_/A VGND VGND VPWR VPWR _2093_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1744_ _1744_/A _1872_/B VGND VGND VPWR VPWR _1968_/A sky130_fd_sc_hd__nand2_2
X_1675_ _2837_/A _2674_/A _3124_/A VGND VGND VPWR VPWR _1675_/X sky130_fd_sc_hd__or3_1
X_3345_ _2417_/Y _2413_/Y _3346_/S VGND VGND VPWR VPWR _3345_/X sky130_fd_sc_hd__mux2_2
X_3276_ _3119_/Y _3117_/Y _3340_/S VGND VGND VPWR VPWR _3276_/X sky130_fd_sc_hd__mux2_1
X_2227_ _2815_/A VGND VGND VPWR VPWR _2359_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2158_ _2158_/A _2812_/A VGND VGND VPWR VPWR _3041_/B sky130_fd_sc_hd__and2_1
X_2089_ _2089_/A _2089_/B VGND VGND VPWR VPWR _2787_/B sky130_fd_sc_hd__nor2_4
XFILLER_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3130_ _2596_/Y _2593_/Y _3346_/S VGND VGND VPWR VPWR _3130_/X sky130_fd_sc_hd__mux2_2
X_3061_ _3099_/C VGND VGND VPWR VPWR _3108_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2012_ _2012_/A VGND VGND VPWR VPWR _2195_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2914_ _2914_/A _2922_/B VGND VGND VPWR VPWR _2914_/X sky130_fd_sc_hd__or2_1
XFILLER_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2845_ _2864_/A _2845_/B VGND VGND VPWR VPWR _2845_/Y sky130_fd_sc_hd__nor2_1
X_2776_ _2776_/A _2776_/B VGND VGND VPWR VPWR _2776_/Y sky130_fd_sc_hd__nor2_1
X_1727_ _1581_/X _2685_/B _1726_/X VGND VGND VPWR VPWR _1727_/Y sky130_fd_sc_hd__o21ai_1
X_1658_ _1670_/A _1658_/B VGND VGND VPWR VPWR _2672_/B sky130_fd_sc_hd__nor2_4
X_1589_ _1589_/A VGND VGND VPWR VPWR _1642_/A sky130_fd_sc_hd__inv_2
X_3328_ _2273_/Y _2851_/B _3351_/S VGND VGND VPWR VPWR _3328_/X sky130_fd_sc_hd__mux2_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3259_ _3059_/Y _3056_/Y _3346_/S VGND VGND VPWR VPWR _3259_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2630_ _2723_/A VGND VGND VPWR VPWR _2630_/X sky130_fd_sc_hd__clkbuf_2
Xoutput217 _3175_/X VGND VGND VPWR VPWR output_thermometer_o[47] sky130_fd_sc_hd__clkbuf_2
X_2561_ _1653_/X _3031_/B _2560_/X VGND VGND VPWR VPWR _2561_/Y sky130_fd_sc_hd__o21ai_1
Xoutput206 _3307_/X VGND VGND VPWR VPWR output_thermometer_o[179] sky130_fd_sc_hd__clkbuf_2
Xoutput239 _3344_/X VGND VGND VPWR VPWR output_thermometer_o[216] sky130_fd_sc_hd__clkbuf_2
X_2492_ _2972_/B VGND VGND VPWR VPWR _2492_/Y sky130_fd_sc_hd__inv_2
Xoutput228 _3155_/X VGND VGND VPWR VPWR output_thermometer_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3113_ _3097_/X _2881_/B _3098_/X _2652_/B _3112_/X VGND VGND VPWR VPWR _3113_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3044_ _3044_/A VGND VGND VPWR VPWR _3044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2828_ _2839_/A _2828_/B VGND VGND VPWR VPWR _2828_/Y sky130_fd_sc_hd__nor2_1
X_2759_ _2759_/A VGND VGND VPWR VPWR _2776_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1992_ _2157_/A VGND VGND VPWR VPWR _1992_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2613_ _2606_/X _2845_/B _2612_/X VGND VGND VPWR VPWR _2613_/Y sky130_fd_sc_hd__o21ai_1
X_2544_ _2788_/A _2990_/B VGND VGND VPWR VPWR _3019_/B sky130_fd_sc_hd__nor2_2
X_2475_ _2509_/B VGND VGND VPWR VPWR _2495_/B sky130_fd_sc_hd__buf_1
XFILLER_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3027_ _3027_/A VGND VGND VPWR VPWR _3041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2260_ _2184_/X _3072_/B _3110_/A VGND VGND VPWR VPWR _2848_/B sky130_fd_sc_hd__o21a_1
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2191_ _2195_/A _2340_/A VGND VGND VPWR VPWR _3048_/B sky130_fd_sc_hd__nor2_2
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1975_ _1951_/X _1970_/A _1961_/X VGND VGND VPWR VPWR _2982_/B sky130_fd_sc_hd__a21oi_4
X_2527_ _2527_/A VGND VGND VPWR VPWR _2527_/X sky130_fd_sc_hd__clkbuf_2
X_2458_ _2946_/B VGND VGND VPWR VPWR _2458_/Y sky130_fd_sc_hd__inv_2
X_2389_ _2184_/A _2387_/B _2142_/A VGND VGND VPWR VPWR _2894_/B sky130_fd_sc_hd__o21a_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1760_ _1884_/A _1884_/B VGND VGND VPWR VPWR _1980_/A sky130_fd_sc_hd__or2_2
X_1691_ _1691_/A VGND VGND VPWR VPWR _2030_/A sky130_fd_sc_hd__clkbuf_2
X_3361_ _2490_/Y _2487_/Y _3365_/S VGND VGND VPWR VPWR _3361_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2312_ _2212_/X _2868_/B _2311_/X VGND VGND VPWR VPWR _2312_/Y sky130_fd_sc_hd__o21ai_1
X_3292_ _1870_/Y _1865_/Y _3357_/S VGND VGND VPWR VPWR _3292_/X sky130_fd_sc_hd__mux2_2
X_2243_ _2400_/A _2243_/B VGND VGND VPWR VPWR _2249_/A sky130_fd_sc_hd__or2_2
X_2174_ _1797_/X _1792_/Y _2171_/X _2173_/X VGND VGND VPWR VPWR _2174_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1958_ _1931_/X _2499_/A _1935_/X VGND VGND VPWR VPWR _1964_/B sky130_fd_sc_hd__o21ai_2
X_1889_ _1938_/A _1889_/B VGND VGND VPWR VPWR _1889_/Y sky130_fd_sc_hd__nor2_1
Xoutput28 _3292_/X VGND VGND VPWR VPWR output_thermometer_o[164] sky130_fd_sc_hd__clkbuf_2
Xoutput17 _3186_/X VGND VGND VPWR VPWR output_thermometer_o[58] sky130_fd_sc_hd__clkbuf_2
Xoutput39 _3330_/X VGND VGND VPWR VPWR output_thermometer_o[202] sky130_fd_sc_hd__clkbuf_2
XFILLER_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2930_ _1769_/C _2920_/X _2921_/X _2694_/B _2929_/X VGND VGND VPWR VPWR _2930_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2861_ _2864_/A _2861_/B VGND VGND VPWR VPWR _2861_/Y sky130_fd_sc_hd__nor2_1
X_2792_ _3022_/A _2792_/B VGND VGND VPWR VPWR _2792_/X sky130_fd_sc_hd__or2_1
X_1812_ _2157_/C VGND VGND VPWR VPWR _2233_/A sky130_fd_sc_hd__buf_2
X_1743_ _3385_/Q _1809_/B _1808_/B VGND VGND VPWR VPWR _1872_/B sky130_fd_sc_hd__o21a_1
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1674_ _3057_/A VGND VGND VPWR VPWR _3124_/A sky130_fd_sc_hd__clkbuf_2
X_3344_ _2412_/Y _2410_/Y _3347_/S VGND VGND VPWR VPWR _3344_/X sky130_fd_sc_hd__mux2_2
X_3275_ _3116_/Y _3114_/Y _3357_/S VGND VGND VPWR VPWR _3275_/X sky130_fd_sc_hd__mux2_1
X_2226_ _2202_/X _2600_/B _2225_/X VGND VGND VPWR VPWR _2226_/Y sky130_fd_sc_hd__o21ai_1
X_2157_ _2157_/A _2157_/B _2157_/C VGND VGND VPWR VPWR _2812_/A sky130_fd_sc_hd__or3_4
X_2088_ _2090_/A _2020_/X _1928_/A _2019_/X _1725_/A VGND VGND VPWR VPWR _3018_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3060_ _3064_/A _3060_/B VGND VGND VPWR VPWR _3060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2011_ _1974_/X _2992_/B _1963_/X _2760_/B _2061_/B VGND VGND VPWR VPWR _2011_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2913_ _2924_/A _2913_/B VGND VGND VPWR VPWR _2913_/Y sky130_fd_sc_hd__nor2_1
X_2844_ _2867_/A VGND VGND VPWR VPWR _2864_/A sky130_fd_sc_hd__clkbuf_2
X_2775_ _2530_/A _2763_/X _3003_/B _2773_/X _2774_/X VGND VGND VPWR VPWR _2775_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1726_ _1708_/X _2421_/A _1622_/X _2916_/B VGND VGND VPWR VPWR _1726_/X sky130_fd_sc_hd__o22a_1
X_1657_ _2193_/A _2889_/A VGND VGND VPWR VPWR _1670_/A sky130_fd_sc_hd__or2_4
X_1588_ _1860_/A VGND VGND VPWR VPWR _1588_/Y sky130_fd_sc_hd__inv_2
X_3327_ _2264_/Y _2254_/Y _3351_/S VGND VGND VPWR VPWR _3327_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3258_ _3055_/Y _3051_/Y _3346_/S VGND VGND VPWR VPWR _3258_/X sky130_fd_sc_hd__mux2_2
X_3189_ _2810_/Y _2808_/Y _3380_/S VGND VGND VPWR VPWR _3189_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2209_ _2202_/X _2593_/B _2208_/X VGND VGND VPWR VPWR _2209_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2560_ _2802_/B _2390_/X _3033_/B _2549_/X VGND VGND VPWR VPWR _2560_/X sky130_fd_sc_hd__o22a_1
Xoutput207 _3245_/X VGND VGND VPWR VPWR output_thermometer_o[117] sky130_fd_sc_hd__clkbuf_2
Xoutput229 _3179_/X VGND VGND VPWR VPWR output_thermometer_o[51] sky130_fd_sc_hd__clkbuf_2
X_2491_ _2491_/A _2495_/B VGND VGND VPWR VPWR _2972_/B sky130_fd_sc_hd__or2_2
Xoutput218 _3275_/X VGND VGND VPWR VPWR output_thermometer_o[147] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3112_ _3124_/A _3112_/B VGND VGND VPWR VPWR _3112_/X sky130_fd_sc_hd__or2_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3043_ _2812_/A _2607_/X _3032_/X _2811_/B _3042_/X VGND VGND VPWR VPWR _3043_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2827_ _2825_/X _3048_/B _1660_/X _2588_/B _2826_/X VGND VGND VPWR VPWR _2827_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2758_ _1996_/B _2743_/X _2989_/B _2753_/X _2788_/B VGND VGND VPWR VPWR _2758_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1709_ _2044_/A VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__clkbuf_2
X_2689_ _2922_/A _2581_/A _2328_/X _2425_/A VGND VGND VPWR VPWR _2689_/X sky130_fd_sc_hd__o22a_1
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1991_ _1991_/A VGND VGND VPWR VPWR _2514_/A sky130_fd_sc_hd__inv_2
X_2612_ _3068_/B _2611_/X _2240_/B _2584_/X VGND VGND VPWR VPWR _2612_/X sky130_fd_sc_hd__o22a_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2543_ _2784_/B _2527_/X _2542_/X VGND VGND VPWR VPWR _2543_/Y sky130_fd_sc_hd__o21ai_1
X_2474_ _2722_/B _2459_/X _2473_/X VGND VGND VPWR VPWR _2474_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3026_ _2795_/A _2920_/X _3015_/X _2794_/B _3025_/X VGND VGND VPWR VPWR _3026_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2190_ _2277_/A VGND VGND VPWR VPWR _2340_/A sky130_fd_sc_hd__buf_2
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1974_ _2087_/A VGND VGND VPWR VPWR _1974_/X sky130_fd_sc_hd__clkbuf_2
X_2526_ _2526_/A _2548_/B VGND VGND VPWR VPWR _2526_/Y sky130_fd_sc_hd__nor2_1
X_2457_ _2457_/A _2471_/B VGND VGND VPWR VPWR _2946_/B sky130_fd_sc_hd__or2_1
XFILLER_68_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2388_ _2388_/A VGND VGND VPWR VPWR _2388_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3009_ _3029_/A _3009_/B VGND VGND VPWR VPWR _3009_/X sky130_fd_sc_hd__or2_1
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1690_ _1722_/A VGND VGND VPWR VPWR _1769_/A sky130_fd_sc_hd__buf_1
X_3360_ _2485_/Y _2482_/Y _3383_/S VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__mux2_2
X_2311_ _2263_/A _3093_/B _2294_/X _2636_/B VGND VGND VPWR VPWR _2311_/X sky130_fd_sc_hd__o22a_1
X_3291_ _1859_/Y _1852_/Y _3383_/S VGND VGND VPWR VPWR _3291_/X sky130_fd_sc_hd__mux2_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2242_ _2242_/A VGND VGND VPWR VPWR _2380_/A sky130_fd_sc_hd__buf_4
X_2173_ _2435_/A VGND VGND VPWR VPWR _2173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1957_ _2298_/B VGND VGND VPWR VPWR _2499_/A sky130_fd_sc_hd__inv_2
X_1888_ _1892_/B VGND VGND VPWR VPWR _1889_/B sky130_fd_sc_hd__inv_2
Xoutput29 _3259_/X VGND VGND VPWR VPWR output_thermometer_o[131] sky130_fd_sc_hd__clkbuf_2
Xoutput18 _3219_/X VGND VGND VPWR VPWR output_thermometer_o[91] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2509_ _2509_/A _2509_/B VGND VGND VPWR VPWR _2986_/B sky130_fd_sc_hd__or2_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2860_ _2857_/X _3083_/B _2833_/X _2625_/B _2859_/X VGND VGND VPWR VPWR _2860_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1811_ _1811_/A VGND VGND VPWR VPWR _2446_/A sky130_fd_sc_hd__inv_2
X_2791_ _2791_/A VGND VGND VPWR VPWR _2791_/X sky130_fd_sc_hd__buf_2
X_1742_ _1735_/X _2688_/B _1741_/X VGND VGND VPWR VPWR _1742_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1673_ _1673_/A VGND VGND VPWR VPWR _2674_/A sky130_fd_sc_hd__inv_2
X_3343_ _2409_/Y _2406_/Y _3346_/S VGND VGND VPWR VPWR _3343_/X sky130_fd_sc_hd__mux2_2
X_3274_ _3113_/Y _3111_/Y _3340_/S VGND VGND VPWR VPWR _3274_/X sky130_fd_sc_hd__mux2_2
X_2225_ _2315_/A _2836_/B _2206_/X _3060_/B VGND VGND VPWR VPWR _2225_/X sky130_fd_sc_hd__o22a_1
X_2156_ _2156_/A _2156_/B VGND VGND VPWR VPWR _2811_/B sky130_fd_sc_hd__nor2_2
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2087_ _2087_/A VGND VGND VPWR VPWR _2087_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2989_ _3003_/A _2989_/B VGND VGND VPWR VPWR _2989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2010_ _2090_/B VGND VGND VPWR VPWR _2061_/B sky130_fd_sc_hd__buf_1
XFILLER_35_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2912_ _1695_/C _2901_/X _2872_/X _2676_/B _2911_/X VGND VGND VPWR VPWR _2912_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2843_ _2087_/X _2605_/B _2840_/X _3065_/B _2842_/X VGND VGND VPWR VPWR _2843_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2774_ _3005_/B _2782_/B VGND VGND VPWR VPWR _2774_/X sky130_fd_sc_hd__or2_1
X_1725_ _1725_/A _1725_/B _1725_/C VGND VGND VPWR VPWR _2916_/B sky130_fd_sc_hd__and3_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1656_ _2168_/B VGND VGND VPWR VPWR _2889_/A sky130_fd_sc_hd__buf_1
X_1587_ _3388_/Q VGND VGND VPWR VPWR _1860_/A sky130_fd_sc_hd__clkbuf_2
X_3326_ _2251_/Y _2241_/Y _3330_/S VGND VGND VPWR VPWR _3326_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3257_ _3050_/Y _3048_/Y _3330_/S VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__mux2_2
X_3188_ _2807_/Y _2805_/Y _3381_/S VGND VGND VPWR VPWR _3188_/X sky130_fd_sc_hd__mux2_1
X_2208_ _2315_/A _2828_/B _2206_/X _3051_/B VGND VGND VPWR VPWR _2208_/X sky130_fd_sc_hd__o22a_1
X_2139_ _2155_/A _3036_/B VGND VGND VPWR VPWR _2139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput208 _3364_/X VGND VGND VPWR VPWR output_thermometer_o[236] sky130_fd_sc_hd__clkbuf_2
Xoutput219 _3158_/X VGND VGND VPWR VPWR output_thermometer_o[30] sky130_fd_sc_hd__clkbuf_2
X_2490_ _2733_/B _2483_/X _2489_/X VGND VGND VPWR VPWR _2490_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3111_ _3126_/A _3111_/B VGND VGND VPWR VPWR _3111_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3042_ _3042_/A _3042_/B VGND VGND VPWR VPWR _3042_/X sky130_fd_sc_hd__or2_1
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2826_ _3049_/B _2854_/B VGND VGND VPWR VPWR _2826_/X sky130_fd_sc_hd__or2_1
X_2757_ _2762_/A _2990_/B VGND VGND VPWR VPWR _2788_/B sky130_fd_sc_hd__or2_1
X_2688_ _2694_/A _2688_/B VGND VGND VPWR VPWR _2688_/Y sky130_fd_sc_hd__nor2_1
X_1708_ _3099_/C VGND VGND VPWR VPWR _1708_/X sky130_fd_sc_hd__clkbuf_2
X_1639_ _2347_/A VGND VGND VPWR VPWR _1639_/X sky130_fd_sc_hd__buf_4
X_3309_ _2072_/Y _2066_/Y _3381_/S VGND VGND VPWR VPWR _3309_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1990_ _1974_/X _2985_/B _1963_/X _2752_/B _1989_/X VGND VGND VPWR VPWR _1990_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_54_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2611_ _2766_/A VGND VGND VPWR VPWR _2611_/X sky130_fd_sc_hd__clkbuf_2
X_2542_ _1653_/A _3014_/B _2075_/B _2531_/X VGND VGND VPWR VPWR _2542_/X sky130_fd_sc_hd__o22a_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2473_ _2454_/X _2955_/B _1889_/B _2464_/X VGND VGND VPWR VPWR _2473_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3025_ _3029_/A _3025_/B VGND VGND VPWR VPWR _3025_/X sky130_fd_sc_hd__or2_1
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2809_ _2809_/A _2849_/A VGND VGND VPWR VPWR _2809_/X sky130_fd_sc_hd__or2_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1973_ _1996_/A _1973_/B VGND VGND VPWR VPWR _1973_/Y sky130_fd_sc_hd__nor2_1
X_2525_ _2765_/B _2506_/X _2524_/X VGND VGND VPWR VPWR _2525_/Y sky130_fd_sc_hd__o21ai_1
X_2456_ _2707_/B _2428_/X _2455_/X VGND VGND VPWR VPWR _2456_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2387_ _3080_/A _2387_/B VGND VGND VPWR VPWR _2388_/A sky130_fd_sc_hd__or2_2
X_3008_ _3024_/A _3008_/B VGND VGND VPWR VPWR _3008_/Y sky130_fd_sc_hd__nor2_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3290_ _1846_/Y _1838_/Y _3354_/S VGND VGND VPWR VPWR _3290_/X sky130_fd_sc_hd__mux2_2
X_2310_ _2310_/A _2344_/A VGND VGND VPWR VPWR _2636_/B sky130_fd_sc_hd__nor2_4
XFILLER_2_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2241_ _3069_/B VGND VGND VPWR VPWR _2241_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2172_ _2578_/A _2582_/B VGND VGND VPWR VPWR _2435_/A sky130_fd_sc_hd__or2_2
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1956_ _1884_/A _1759_/A _1588_/Y VGND VGND VPWR VPWR _2298_/B sky130_fd_sc_hd__o21ai_4
X_1887_ _1871_/X _2471_/A _1875_/X VGND VGND VPWR VPWR _1892_/B sky130_fd_sc_hd__o21ai_2
Xoutput19 _3192_/X VGND VGND VPWR VPWR output_thermometer_o[64] sky130_fd_sc_hd__clkbuf_2
X_2508_ _2749_/B _2506_/X _2507_/X VGND VGND VPWR VPWR _2508_/Y sky130_fd_sc_hd__o21ai_1
X_2439_ _2549_/A VGND VGND VPWR VPWR _2803_/B sky130_fd_sc_hd__clkbuf_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1810_ _2067_/A _2012_/A VGND VGND VPWR VPWR _1811_/A sky130_fd_sc_hd__or2_2
XFILLER_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2790_ _2794_/A _2790_/B VGND VGND VPWR VPWR _2790_/Y sky130_fd_sc_hd__nor2_1
X_1741_ _1708_/X _2425_/A _1622_/X _2919_/B VGND VGND VPWR VPWR _1741_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1672_ _2841_/A VGND VGND VPWR VPWR _2837_/A sky130_fd_sc_hd__clkbuf_2
X_3342_ _2405_/Y _2399_/Y _3342_/S VGND VGND VPWR VPWR _3342_/X sky130_fd_sc_hd__mux2_2
X_3273_ _3109_/Y _3107_/Y _3340_/S VGND VGND VPWR VPWR _3273_/X sky130_fd_sc_hd__mux2_1
X_2224_ _2224_/A VGND VGND VPWR VPWR _3060_/B sky130_fd_sc_hd__inv_2
X_2155_ _2155_/A _3042_/B VGND VGND VPWR VPWR _2155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2086_ _2109_/A _2086_/B VGND VGND VPWR VPWR _2086_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2988_ _3027_/A VGND VGND VPWR VPWR _3003_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1939_ _1890_/X _1934_/A _1900_/X VGND VGND VPWR VPWR _2971_/B sky130_fd_sc_hd__a21oi_4
XFILLER_17_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2911_ _2911_/A _2922_/B VGND VGND VPWR VPWR _2911_/X sky130_fd_sc_hd__or2_1
X_2842_ _2887_/A _3064_/B _2879_/C VGND VGND VPWR VPWR _2842_/X sky130_fd_sc_hd__or3_2
X_2773_ _2791_/A VGND VGND VPWR VPWR _2773_/X sky130_fd_sc_hd__clkbuf_2
X_1724_ _2185_/A _1725_/C VGND VGND VPWR VPWR _2421_/A sky130_fd_sc_hd__or2_2
XFILLER_7_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1655_ _1839_/A VGND VGND VPWR VPWR _2193_/A sky130_fd_sc_hd__buf_2
X_1586_ _2257_/A VGND VGND VPWR VPWR _2090_/A sky130_fd_sc_hd__inv_2
X_3325_ _2238_/Y _2230_/Y _3342_/S VGND VGND VPWR VPWR _3325_/X sky130_fd_sc_hd__mux2_2
X_3256_ _3046_/Y _1779_/A _3346_/S VGND VGND VPWR VPWR _3256_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2207_ _2207_/A _2340_/A VGND VGND VPWR VPWR _3051_/B sky130_fd_sc_hd__nor2_2
X_3187_ _2804_/Y _2802_/Y _3380_/S VGND VGND VPWR VPWR _3187_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2138_ _2140_/B VGND VGND VPWR VPWR _3036_/B sky130_fd_sc_hd__inv_2
X_2069_ _1951_/X _2386_/B _1900_/A VGND VGND VPWR VPWR _3011_/B sky130_fd_sc_hd__a21oi_4
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput209 _3242_/X VGND VGND VPWR VPWR output_thermometer_o[114] sky130_fd_sc_hd__clkbuf_2
X_3110_ _3110_/A VGND VGND VPWR VPWR _3126_/A sky130_fd_sc_hd__buf_2
X_3041_ _3041_/A _3041_/B VGND VGND VPWR VPWR _3041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2825_ _2857_/A VGND VGND VPWR VPWR _2825_/X sky130_fd_sc_hd__buf_2
X_2756_ _2756_/A _2756_/B VGND VGND VPWR VPWR _2756_/Y sky130_fd_sc_hd__nor2_1
X_2687_ _2916_/B _2682_/X _2686_/X VGND VGND VPWR VPWR _2687_/Y sky130_fd_sc_hd__o21ai_1
X_1707_ _2089_/A _1707_/B VGND VGND VPWR VPWR _2681_/B sky130_fd_sc_hd__nor2_2
X_1638_ _2568_/A VGND VGND VPWR VPWR _2410_/A sky130_fd_sc_hd__clkbuf_2
X_1569_ _3389_/Q _3388_/Q _3390_/Q VGND VGND VPWR VPWR _2329_/B sky130_fd_sc_hd__or3_4
XFILLER_48_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3308_ _2062_/Y _2056_/Y _3374_/S VGND VGND VPWR VPWR _3308_/X sky130_fd_sc_hd__mux2_4
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3239_ _2991_/Y _2989_/Y _3370_/S VGND VGND VPWR VPWR _3239_/X sky130_fd_sc_hd__mux2_2
XFILLER_54_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2610_ _2610_/A _2610_/B VGND VGND VPWR VPWR _2610_/Y sky130_fd_sc_hd__nor2_1
X_2541_ _2785_/A _2785_/B VGND VGND VPWR VPWR _3016_/B sky130_fd_sc_hd__nor2_1
X_2472_ _2956_/B VGND VGND VPWR VPWR _2472_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3024_ _3024_/A _3024_/B VGND VGND VPWR VPWR _3024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2808_ _2811_/A _2808_/B VGND VGND VPWR VPWR _2808_/Y sky130_fd_sc_hd__nor2_1
X_2739_ _1938_/B _2723_/X _2971_/B _2734_/X _2738_/X VGND VGND VPWR VPWR _2739_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1972_ _1977_/B VGND VGND VPWR VPWR _1973_/B sky130_fd_sc_hd__inv_2
X_2524_ _2523_/X _2996_/B _2998_/B _2511_/X VGND VGND VPWR VPWR _2524_/X sky130_fd_sc_hd__o22a_1
X_2455_ _2454_/X _2938_/B _1838_/B _2436_/X VGND VGND VPWR VPWR _2455_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2386_ _2386_/A _2386_/B VGND VGND VPWR VPWR _2387_/B sky130_fd_sc_hd__nor2_1
XFILLER_56_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3007_ _3027_/A VGND VGND VPWR VPWR _3024_/A sky130_fd_sc_hd__clkbuf_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2240_ _2359_/A _2240_/B VGND VGND VPWR VPWR _3069_/B sky130_fd_sc_hd__or2_2
X_2171_ _2171_/A VGND VGND VPWR VPWR _2171_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1955_ _1913_/X _2974_/B _1902_/X _2741_/B _1954_/X VGND VGND VPWR VPWR _1955_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1886_ _2243_/B VGND VGND VPWR VPWR _2471_/A sky130_fd_sc_hd__inv_2
X_2507_ _2501_/X _2982_/B _1973_/B _2488_/X VGND VGND VPWR VPWR _2507_/X sky130_fd_sc_hd__o22a_1
X_2438_ _2694_/B _2428_/X _2437_/X VGND VGND VPWR VPWR _2438_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2369_ _3115_/B VGND VGND VPWR VPWR _2369_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1740_ _1769_/A _1769_/B _1740_/C VGND VGND VPWR VPWR _2919_/B sky130_fd_sc_hd__and3_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1671_ _1722_/A VGND VGND VPWR VPWR _2841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3341_ _2396_/Y _2388_/Y _3382_/S VGND VGND VPWR VPWR _3341_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3272_ _3106_/Y _3104_/Y _3357_/S VGND VGND VPWR VPWR _3272_/X sky130_fd_sc_hd__mux2_1
X_2223_ _1631_/B _2219_/B _1779_/A VGND VGND VPWR VPWR _2836_/B sky130_fd_sc_hd__a21oi_4
XFILLER_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2154_ _2156_/B VGND VGND VPWR VPWR _3042_/B sky130_fd_sc_hd__inv_2
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2085_ _2089_/B VGND VGND VPWR VPWR _2086_/B sky130_fd_sc_hd__inv_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2987_ _2978_/X _1985_/B _2979_/X _2752_/B _2986_/X VGND VGND VPWR VPWR _2987_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1938_ _1938_/A _1938_/B VGND VGND VPWR VPWR _1938_/Y sky130_fd_sc_hd__nor2_1
X_1869_ _1917_/A _2462_/A _1893_/C VGND VGND VPWR VPWR _1869_/X sky130_fd_sc_hd__or3_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2910_ _2924_/A _2910_/B VGND VGND VPWR VPWR _2910_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2841_ _2841_/A VGND VGND VPWR VPWR _2887_/A sky130_fd_sc_hd__buf_1
X_2772_ _2776_/A _2772_/B VGND VGND VPWR VPWR _2772_/Y sky130_fd_sc_hd__nor2_1
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _2386_/A _1718_/B _1709_/X VGND VGND VPWR VPWR _1725_/C sky130_fd_sc_hd__o21ai_1
X_1654_ _2578_/A VGND VGND VPWR VPWR _1839_/A sky130_fd_sc_hd__inv_2
X_1585_ _3387_/Q _1641_/B VGND VGND VPWR VPWR _2257_/A sky130_fd_sc_hd__or2_2
X_3324_ _2226_/Y _2220_/Y _3346_/S VGND VGND VPWR VPWR _3324_/X sky130_fd_sc_hd__mux2_2
X_3255_ _3045_/X _3044_/X _3354_/S VGND VGND VPWR VPWR _3255_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2206_ _2549_/A VGND VGND VPWR VPWR _2206_/X sky130_fd_sc_hd__buf_2
X_3186_ _2801_/Y _2798_/Y _3380_/S VGND VGND VPWR VPWR _3186_/X sky130_fd_sc_hd__mux2_1
X_2137_ _1988_/A _2141_/B _2291_/A VGND VGND VPWR VPWR _2140_/B sky130_fd_sc_hd__o21ai_4
XFILLER_66_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2068_ _2537_/A VGND VGND VPWR VPWR _2386_/B sky130_fd_sc_hd__inv_2
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3040_ _2809_/A _2607_/X _3032_/X _2808_/B _3039_/X VGND VGND VPWR VPWR _3040_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2824_ _2939_/A VGND VGND VPWR VPWR _2857_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2755_ _1985_/B _2743_/X _2985_/B _2753_/X _2754_/X VGND VGND VPWR VPWR _2755_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2686_ _2917_/A _2581_/A _2393_/X _2421_/A VGND VGND VPWR VPWR _2686_/X sky130_fd_sc_hd__o22a_1
X_1706_ _2410_/A _2914_/A VGND VGND VPWR VPWR _1706_/Y sky130_fd_sc_hd__nor2_1
X_1637_ _2898_/A VGND VGND VPWR VPWR _2568_/A sky130_fd_sc_hd__buf_2
X_3307_ _2053_/Y _2047_/Y _3374_/S VGND VGND VPWR VPWR _3307_/X sky130_fd_sc_hd__mux2_2
X_1568_ _1589_/A VGND VGND VPWR VPWR _1570_/A sky130_fd_sc_hd__clkbuf_2
X_3238_ _2987_/Y _2985_/Y _3370_/S VGND VGND VPWR VPWR _3238_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3169_ _2736_/Y _2733_/Y _3365_/S VGND VGND VPWR VPWR _3169_/X sky130_fd_sc_hd__mux2_4
XFILLER_64_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2540_ _2781_/B _2527_/X _2539_/X VGND VGND VPWR VPWR _2540_/Y sky130_fd_sc_hd__o21ai_1
X_2471_ _2471_/A _2471_/B VGND VGND VPWR VPWR _2956_/B sky130_fd_sc_hd__or2_1
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk_i clk_i VGND VGND VPWR VPWR clkbuf_0_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_3023_ _2857_/A _2095_/B _3015_/X _2790_/B _3022_/X VGND VGND VPWR VPWR _3023_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_36_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_clk_i clkbuf_0_clk_i/X VGND VGND VPWR VPWR _3408_/CLK sky130_fd_sc_hd__clkbuf_1
X_2807_ _3036_/B _2799_/X _3035_/B _2791_/X _2806_/X VGND VGND VPWR VPWR _2807_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2738_ _2744_/A _2972_/B VGND VGND VPWR VPWR _2738_/X sky130_fd_sc_hd__or2_1
X_2669_ _2676_/A _2669_/B VGND VGND VPWR VPWR _2669_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1971_ _1931_/X _2504_/A _1935_/X VGND VGND VPWR VPWR _1977_/B sky130_fd_sc_hd__o21ai_2
XFILLER_60_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2523_ _2523_/A VGND VGND VPWR VPWR _2523_/X sky130_fd_sc_hd__clkbuf_2
X_2454_ _2478_/A VGND VGND VPWR VPWR _2454_/X sky130_fd_sc_hd__clkbuf_2
X_2385_ _2351_/X _2659_/B _2384_/X VGND VGND VPWR VPWR _2385_/Y sky130_fd_sc_hd__o21ai_1
Xinput1 rst_ni VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_6
X_3006_ _2530_/A _2994_/X _2997_/X _2772_/B _3005_/X VGND VGND VPWR VPWR _3006_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2170_ _2390_/A VGND VGND VPWR VPWR _2171_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1954_ _1978_/A _2495_/A _1954_/C VGND VGND VPWR VPWR _1954_/X sky130_fd_sc_hd__or3_2
X_1885_ _1907_/A _2076_/B VGND VGND VPWR VPWR _2243_/B sky130_fd_sc_hd__or2_4
X_2506_ _2527_/A VGND VGND VPWR VPWR _2506_/X sky130_fd_sc_hd__clkbuf_2
X_2437_ _2422_/X _2928_/B _2929_/A _2436_/X VGND VGND VPWR VPWR _2437_/X sky130_fd_sc_hd__o22a_1
X_2368_ _2398_/A _2657_/A VGND VGND VPWR VPWR _3115_/B sky130_fd_sc_hd__or2_2
X_2299_ _2359_/A _2299_/B VGND VGND VPWR VPWR _3091_/B sky130_fd_sc_hd__or2_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput190 _3306_/X VGND VGND VPWR VPWR output_thermometer_o[178] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1670_ _1670_/A _1673_/A VGND VGND VPWR VPWR _2905_/B sky130_fd_sc_hd__nor2_4
X_3340_ _2385_/Y _2378_/Y _3340_/S VGND VGND VPWR VPWR _3340_/X sky130_fd_sc_hd__mux2_1
X_3271_ _3103_/X _3101_/Y _3354_/S VGND VGND VPWR VPWR _3271_/X sky130_fd_sc_hd__mux2_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2222_ _2232_/A _2224_/A VGND VGND VPWR VPWR _2600_/B sky130_fd_sc_hd__nor2_2
X_2153_ _2042_/A _2318_/A _1684_/A _1605_/B VGND VGND VPWR VPWR _2156_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2084_ _2257_/A _2005_/X _2397_/A _2014_/X VGND VGND VPWR VPWR _2089_/B sky130_fd_sc_hd__a31o_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2986_ _2990_/A _2986_/B VGND VGND VPWR VPWR _2986_/X sky130_fd_sc_hd__or2_1
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1937_ _1940_/B VGND VGND VPWR VPWR _1938_/B sky130_fd_sc_hd__inv_2
X_1868_ _1928_/A VGND VGND VPWR VPWR _1917_/A sky130_fd_sc_hd__buf_1
X_1799_ _1799_/A VGND VGND VPWR VPWR _1799_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2840_ _2936_/A VGND VGND VPWR VPWR _2840_/X sky130_fd_sc_hd__clkbuf_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _2526_/A _2763_/X _3000_/B _2753_/X _2770_/X VGND VGND VPWR VPWR _2771_/Y
+ sky130_fd_sc_hd__o221ai_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1722_ _1722_/A VGND VGND VPWR VPWR _2185_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1653_ _1653_/A VGND VGND VPWR VPWR _1653_/X sky130_fd_sc_hd__clkbuf_2
X_1584_ _1584_/A VGND VGND VPWR VPWR _1641_/B sky130_fd_sc_hd__inv_2
X_3323_ _2217_/Y _2211_/Y _3346_/S VGND VGND VPWR VPWR _3323_/X sky130_fd_sc_hd__mux2_2
X_3254_ _3043_/Y _3041_/Y _3382_/S VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__mux2_2
X_2205_ _1631_/B _2199_/B _1779_/A VGND VGND VPWR VPWR _2828_/B sky130_fd_sc_hd__a21oi_4
X_3185_ _2796_/Y _2794_/Y _3381_/S VGND VGND VPWR VPWR _3185_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2136_ _2131_/X _2802_/B _2135_/X VGND VGND VPWR VPWR _2136_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2067_ _2067_/A _2067_/B VGND VGND VPWR VPWR _2537_/A sky130_fd_sc_hd__nand2_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2969_ _2959_/X _1925_/B _2960_/X _2733_/B _2968_/X VGND VGND VPWR VPWR _2969_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2823_ _2839_/A _2823_/B VGND VGND VPWR VPWR _2823_/Y sky130_fd_sc_hd__nor2_1
X_2754_ _2785_/C _2986_/B VGND VGND VPWR VPWR _2754_/X sky130_fd_sc_hd__or2_1
X_1705_ _1707_/B VGND VGND VPWR VPWR _2914_/A sky130_fd_sc_hd__inv_2
X_2685_ _2694_/A _2685_/B VGND VGND VPWR VPWR _2685_/Y sky130_fd_sc_hd__nor2_1
X_1636_ _2234_/A VGND VGND VPWR VPWR _2898_/A sky130_fd_sc_hd__clkbuf_2
X_1567_ _3387_/Q _1584_/A VGND VGND VPWR VPWR _1589_/A sky130_fd_sc_hd__or2_1
X_3306_ _2041_/Y _2033_/Y _3374_/S VGND VGND VPWR VPWR _3306_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3237_ _2984_/Y _2982_/Y _3370_/S VGND VGND VPWR VPWR _3237_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3168_ _2732_/Y _2730_/Y _3383_/S VGND VGND VPWR VPWR _3168_/X sky130_fd_sc_hd__mux2_1
X_2119_ _2042_/X _2286_/A _1684_/A _2044_/X VGND VGND VPWR VPWR _2122_/B sky130_fd_sc_hd__a31o_2
XFILLER_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3099_ _3099_/A _3099_/B _3099_/C VGND VGND VPWR VPWR _3099_/X sky130_fd_sc_hd__or3_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2470_ _2718_/B _2459_/X _2469_/X VGND VGND VPWR VPWR _2470_/Y sky130_fd_sc_hd__o21ai_1
X_3022_ _3022_/A _3022_/B VGND VGND VPWR VPWR _3022_/X sky130_fd_sc_hd__or2_1
X_2806_ _2806_/A _2849_/A VGND VGND VPWR VPWR _2806_/X sky130_fd_sc_hd__or2_1
X_2737_ _2737_/A _2737_/B VGND VGND VPWR VPWR _2737_/Y sky130_fd_sc_hd__nor2_1
X_2668_ _2606_/X _2897_/B _2667_/X VGND VGND VPWR VPWR _2668_/Y sky130_fd_sc_hd__o21ai_1
X_1619_ _2582_/B VGND VGND VPWR VPWR _2762_/A sky130_fd_sc_hd__clkbuf_2
X_2599_ _3056_/B _2581_/X _2594_/X _2831_/B _2598_/X VGND VGND VPWR VPWR _2599_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_27_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1970_ _1970_/A VGND VGND VPWR VPWR _2504_/A sky130_fd_sc_hd__inv_2
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2522_ _2522_/A _2548_/B VGND VGND VPWR VPWR _2522_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2453_ _2943_/B VGND VGND VPWR VPWR _2453_/Y sky130_fd_sc_hd__inv_2
X_2384_ _2381_/X _2891_/B _2248_/X _3117_/B VGND VGND VPWR VPWR _2384_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 randomise_en_i VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3005_ _3029_/A _3005_/B VGND VGND VPWR VPWR _3005_/X sky130_fd_sc_hd__or2_1
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1953_ _1964_/A _1953_/B VGND VGND VPWR VPWR _2741_/B sky130_fd_sc_hd__nor2_2
X_1884_ _1884_/A _1884_/B VGND VGND VPWR VPWR _2076_/B sky130_fd_sc_hd__nand2_2
X_2505_ _2983_/B VGND VGND VPWR VPWR _2505_/Y sky130_fd_sc_hd__inv_2
X_2436_ _2531_/A VGND VGND VPWR VPWR _2436_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2367_ _2347_/X _2049_/A _2009_/B VGND VGND VPWR VPWR _2657_/A sky130_fd_sc_hd__o21a_1
X_2298_ _2386_/A _2298_/B VGND VGND VPWR VPWR _2299_/B sky130_fd_sc_hd__nor2_2
XFILLER_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput180 _3229_/X VGND VGND VPWR VPWR output_thermometer_o[101] sky130_fd_sc_hd__clkbuf_2
Xoutput191 _3214_/X VGND VGND VPWR VPWR output_thermometer_o[86] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3270_ _3100_/Y _3096_/Y _3340_/S VGND VGND VPWR VPWR _3270_/X sky130_fd_sc_hd__mux2_1
X_2221_ _2400_/A _2221_/B VGND VGND VPWR VPWR _2224_/A sky130_fd_sc_hd__or2_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2152_ _2131_/X _2808_/B _2151_/X VGND VGND VPWR VPWR _2152_/Y sky130_fd_sc_hd__o21ai_1
X_2083_ _2034_/X _3014_/B _2080_/X _2784_/B _2082_/X VGND VGND VPWR VPWR _2083_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2985_ _2985_/A _2985_/B VGND VGND VPWR VPWR _2985_/Y sky130_fd_sc_hd__nor2_1
X_1936_ _1931_/X _2491_/A _1935_/X VGND VGND VPWR VPWR _1940_/B sky130_fd_sc_hd__o21ai_2
X_1867_ _1903_/A _1867_/B VGND VGND VPWR VPWR _2714_/B sky130_fd_sc_hd__nor2_4
X_1798_ _1624_/B _2391_/A _2391_/C VGND VGND VPWR VPWR _1799_/A sky130_fd_sc_hd__o21ai_2
X_2419_ _2381_/X _2913_/B _2914_/A _2415_/X VGND VGND VPWR VPWR _2419_/X sky130_fd_sc_hd__o22a_1
X_3399_ _3404_/CLK _3399_/D input1/X VGND VGND VPWR VPWR _3400_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_37_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _3001_/B _2782_/B VGND VGND VPWR VPWR _2770_/X sky130_fd_sc_hd__or2_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _2089_/A _1721_/B VGND VGND VPWR VPWR _2685_/B sky130_fd_sc_hd__nor2_2
X_1652_ _2523_/A VGND VGND VPWR VPWR _1653_/A sky130_fd_sc_hd__clkbuf_2
X_1583_ _2333_/A VGND VGND VPWR VPWR _2401_/A sky130_fd_sc_hd__clkbuf_4
X_3322_ _2209_/Y _2200_/Y _3346_/S VGND VGND VPWR VPWR _3322_/X sky130_fd_sc_hd__mux2_2
X_3253_ _3040_/Y _3038_/Y _3380_/S VGND VGND VPWR VPWR _3253_/X sky130_fd_sc_hd__mux2_1
X_3184_ _2793_/Y _2790_/Y _3374_/S VGND VGND VPWR VPWR _3184_/X sky130_fd_sc_hd__mux2_2
X_2204_ _3098_/A VGND VGND VPWR VPWR _2315_/A sky130_fd_sc_hd__clkbuf_2
X_2135_ _1755_/X _3031_/B _2133_/B _1802_/X VGND VGND VPWR VPWR _2135_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2066_ _2109_/A _3012_/B VGND VGND VPWR VPWR _2066_/Y sky130_fd_sc_hd__nor2_1
X_2968_ _2975_/A _2968_/B VGND VGND VPWR VPWR _2968_/X sky130_fd_sc_hd__or2_1
X_1919_ _2076_/A VGND VGND VPWR VPWR _1981_/A sky130_fd_sc_hd__buf_1
X_2899_ _2882_/X _2666_/B _2331_/X _3124_/B _2898_/X VGND VGND VPWR VPWR _2899_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_1_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2822_ _2867_/A VGND VGND VPWR VPWR _2839_/A sky130_fd_sc_hd__clkbuf_2
X_2753_ _2791_/A VGND VGND VPWR VPWR _2753_/X sky130_fd_sc_hd__clkbuf_2
X_1704_ _1763_/A _1704_/B _1747_/C VGND VGND VPWR VPWR _1707_/B sky130_fd_sc_hd__or3_4
X_2684_ _2913_/B _2682_/X _2683_/X VGND VGND VPWR VPWR _2684_/Y sky130_fd_sc_hd__o21ai_1
X_1635_ _1722_/A VGND VGND VPWR VPWR _2234_/A sky130_fd_sc_hd__clkbuf_2
X_1566_ _1566_/A _1847_/A VGND VGND VPWR VPWR _1584_/A sky130_fd_sc_hd__nand2_2
X_3305_ _2028_/Y _2017_/Y _3374_/S VGND VGND VPWR VPWR _3305_/X sky130_fd_sc_hd__mux2_1
X_3236_ _2981_/Y _2977_/Y _3365_/S VGND VGND VPWR VPWR _3236_/X sky130_fd_sc_hd__mux2_2
X_3167_ _2729_/Y _2726_/Y _3383_/S VGND VGND VPWR VPWR _3167_/X sky130_fd_sc_hd__mux2_4
X_2118_ _3047_/A VGND VGND VPWR VPWR _2155_/A sky130_fd_sc_hd__clkbuf_2
X_3098_ _3098_/A VGND VGND VPWR VPWR _3098_/X sky130_fd_sc_hd__clkbuf_2
X_2049_ _2049_/A VGND VGND VPWR VPWR _2530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3021_ _3021_/A VGND VGND VPWR VPWR _3021_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2805_ _2811_/A _2805_/B VGND VGND VPWR VPWR _2805_/Y sky130_fd_sc_hd__nor2_1
X_2736_ _1925_/B _2723_/X _2967_/B _2734_/X _2735_/X VGND VGND VPWR VPWR _2736_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2667_ _3123_/B _2611_/X _2398_/B _2618_/B VGND VGND VPWR VPWR _2667_/X sky130_fd_sc_hd__o22a_1
X_1618_ _1618_/A _2577_/B VGND VGND VPWR VPWR _2582_/B sky130_fd_sc_hd__or2_1
X_2598_ _3058_/B _2618_/B VGND VGND VPWR VPWR _2598_/X sky130_fd_sc_hd__or2_1
X_3219_ _2918_/Y _2916_/Y _3347_/S VGND VGND VPWR VPWR _3219_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2521_ _2993_/B VGND VGND VPWR VPWR _2548_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2452_ _2452_/A _2471_/B VGND VGND VPWR VPWR _2943_/B sky130_fd_sc_hd__or2_1
XFILLER_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2383_ _2383_/A VGND VGND VPWR VPWR _3117_/B sky130_fd_sc_hd__inv_2
XFILLER_68_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3004_ _3004_/A VGND VGND VPWR VPWR _3029_/A sky130_fd_sc_hd__buf_1
Xinput3 input_binary_i[0] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2719_ _2724_/A _2953_/B VGND VGND VPWR VPWR _2719_/X sky130_fd_sc_hd__or2_1
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ _1951_/X _1947_/A _1900_/X VGND VGND VPWR VPWR _2974_/B sky130_fd_sc_hd__a21oi_4
X_1883_ _2568_/A VGND VGND VPWR VPWR _1938_/A sky130_fd_sc_hd__clkbuf_2
X_2504_ _2504_/A _2509_/B VGND VGND VPWR VPWR _2983_/B sky130_fd_sc_hd__or2_1
X_2435_ _2435_/A VGND VGND VPWR VPWR _2531_/A sky130_fd_sc_hd__buf_2
X_2366_ _2351_/X _2652_/B _2365_/X VGND VGND VPWR VPWR _2366_/Y sky130_fd_sc_hd__o21ai_1
X_2297_ _2212_/X _2861_/B _2296_/X VGND VGND VPWR VPWR _2297_/Y sky130_fd_sc_hd__o21ai_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput170 _3296_/X VGND VGND VPWR VPWR output_thermometer_o[168] sky130_fd_sc_hd__clkbuf_2
Xoutput192 _3316_/X VGND VGND VPWR VPWR output_thermometer_o[188] sky130_fd_sc_hd__clkbuf_2
Xoutput181 _3239_/X VGND VGND VPWR VPWR output_thermometer_o[111] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2220_ _3062_/B VGND VGND VPWR VPWR _2220_/Y sky130_fd_sc_hd__inv_2
X_2151_ _1818_/A _3038_/B _2149_/B _1802_/A VGND VGND VPWR VPWR _2151_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2082_ _2082_/A _2785_/A _2082_/C VGND VGND VPWR VPWR _2082_/X sky130_fd_sc_hd__or3_1
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2984_ _2978_/X _1973_/B _2979_/X _2749_/B _2983_/X VGND VGND VPWR VPWR _2984_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_61_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1935_ _2233_/A VGND VGND VPWR VPWR _1935_/X sky130_fd_sc_hd__buf_2
X_1866_ _1820_/X _2221_/B _1840_/X VGND VGND VPWR VPWR _2948_/B sky130_fd_sc_hd__a21oi_4
X_1797_ _2936_/A VGND VGND VPWR VPWR _1797_/X sky130_fd_sc_hd__buf_2
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2418_ _2418_/A VGND VGND VPWR VPWR _2418_/Y sky130_fd_sc_hd__inv_2
X_3398_ _3404_/CLK _3398_/D input1/X VGND VGND VPWR VPWR _3399_/D sky130_fd_sc_hd__dfrtp_1
X_2349_ _2359_/A _2650_/A VGND VGND VPWR VPWR _3108_/B sky130_fd_sc_hd__or2_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1720_ _2410_/A _2917_/A VGND VGND VPWR VPWR _1720_/Y sky130_fd_sc_hd__nor2_1
X_1651_ _2410_/A _2907_/A VGND VGND VPWR VPWR _1651_/Y sky130_fd_sc_hd__nor2_1
X_1582_ _3391_/Q VGND VGND VPWR VPWR _2333_/A sky130_fd_sc_hd__buf_1
X_3321_ _2197_/Y _2182_/Y _3346_/S VGND VGND VPWR VPWR _3321_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3252_ _3037_/Y _3035_/Y _3381_/S VGND VGND VPWR VPWR _3252_/X sky130_fd_sc_hd__mux2_1
X_3183_ _2789_/Y _2787_/Y _3374_/S VGND VGND VPWR VPWR _3183_/X sky130_fd_sc_hd__mux2_2
X_2203_ _2207_/A _2286_/B VGND VGND VPWR VPWR _2593_/B sky130_fd_sc_hd__nor2_2
X_2134_ _2158_/A _2803_/A VGND VGND VPWR VPWR _3031_/B sky130_fd_sc_hd__and2_1
X_2065_ _2070_/B VGND VGND VPWR VPWR _3012_/B sky130_fd_sc_hd__inv_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2967_ _2967_/A _2967_/B VGND VGND VPWR VPWR _2967_/Y sky130_fd_sc_hd__nor2_1
X_2898_ _2898_/A _3123_/B _3049_/C VGND VGND VPWR VPWR _2898_/X sky130_fd_sc_hd__or3_2
X_1918_ _1913_/X _2964_/B _1902_/X _2730_/B _1917_/X VGND VGND VPWR VPWR _1918_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1849_ _1849_/A VGND VGND VPWR VPWR _2457_/A sky130_fd_sc_hd__inv_2
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2821_ _2854_/B _2821_/B VGND VGND VPWR VPWR _2821_/Y sky130_fd_sc_hd__nand2_1
X_2752_ _2756_/A _2752_/B VGND VGND VPWR VPWR _2752_/Y sky130_fd_sc_hd__nor2_1
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1703_ _2124_/B VGND VGND VPWR VPWR _1704_/B sky130_fd_sc_hd__inv_2
X_2683_ _2914_/A _2611_/X _2393_/X _2418_/A VGND VGND VPWR VPWR _2683_/X sky130_fd_sc_hd__o22a_1
X_1634_ _1581_/X _2669_/B _1633_/X VGND VGND VPWR VPWR _1634_/Y sky130_fd_sc_hd__o21ai_1
X_1565_ _3385_/Q _3384_/Q VGND VGND VPWR VPWR _1847_/A sky130_fd_sc_hd__nor2_8
X_3304_ _2011_/Y _2004_/Y _3374_/S VGND VGND VPWR VPWR _3304_/X sky130_fd_sc_hd__mux2_4
X_3235_ _2976_/Y _2974_/Y _3365_/S VGND VGND VPWR VPWR _3235_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3166_ _2725_/Y _2722_/Y _3383_/S VGND VGND VPWR VPWR _3166_/X sky130_fd_sc_hd__mux2_1
X_2117_ _1735_/X _2794_/B _2116_/X VGND VGND VPWR VPWR _2117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3097_ _3097_/A VGND VGND VPWR VPWR _3097_/X sky130_fd_sc_hd__clkbuf_2
X_2048_ _2215_/A VGND VGND VPWR VPWR _2049_/A sky130_fd_sc_hd__inv_2
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3020_ _2857_/A _2086_/B _3015_/X _2787_/B _3019_/Y VGND VGND VPWR VPWR _3020_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2804_ _3033_/B _2799_/X _3031_/B _2791_/X _2803_/X VGND VGND VPWR VPWR _2804_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2735_ _2744_/A _2968_/B VGND VGND VPWR VPWR _2735_/X sky130_fd_sc_hd__or2_1
X_2666_ _2676_/A _2666_/B VGND VGND VPWR VPWR _2666_/Y sky130_fd_sc_hd__nor2_1
X_1617_ _3102_/A VGND VGND VPWR VPWR _2577_/B sky130_fd_sc_hd__inv_2
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2597_ _2610_/A _2597_/B VGND VGND VPWR VPWR _2597_/Y sky130_fd_sc_hd__nor2_1
X_3218_ _2915_/Y _2913_/Y _3347_/S VGND VGND VPWR VPWR _3218_/X sky130_fd_sc_hd__mux2_2
X_3149_ _2665_/Y _2663_/Y _3382_/S VGND VGND VPWR VPWR _3149_/X sky130_fd_sc_hd__mux2_2
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2520_ _2760_/B _2506_/X _2519_/X VGND VGND VPWR VPWR _2520_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2451_ _2509_/B VGND VGND VPWR VPWR _2471_/B sky130_fd_sc_hd__buf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2382_ _2233_/X _2660_/A _2234_/X VGND VGND VPWR VPWR _2891_/B sky130_fd_sc_hd__o21a_1
XFILLER_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3003_ _3003_/A _3003_/B VGND VGND VPWR VPWR _3003_/Y sky130_fd_sc_hd__nor2_1
Xinput4 input_binary_i[1] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2718_ _2718_/A _2718_/B VGND VGND VPWR VPWR _2718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2649_ _2659_/A _2649_/B VGND VGND VPWR VPWR _2649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1951_ _1951_/A VGND VGND VPWR VPWR _1951_/X sky130_fd_sc_hd__buf_4
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1882_ _1854_/X _2952_/B _1842_/X _2718_/B _1881_/X VGND VGND VPWR VPWR _1882_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2503_ _2746_/B _2483_/X _2502_/X VGND VGND VPWR VPWR _2503_/Y sky130_fd_sc_hd__o21ai_1
X_2434_ _2434_/A VGND VGND VPWR VPWR _2434_/Y sky130_fd_sc_hd__inv_2
X_2365_ _2246_/X _2881_/B _2248_/X _3111_/B VGND VGND VPWR VPWR _2365_/X sky130_fd_sc_hd__o22a_1
X_2296_ _2263_/A _3087_/B _2294_/X _2629_/B VGND VGND VPWR VPWR _2296_/X sky130_fd_sc_hd__o22a_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput160 _3181_/X VGND VGND VPWR VPWR output_thermometer_o[53] sky130_fd_sc_hd__clkbuf_2
Xoutput193 _3328_/X VGND VGND VPWR VPWR output_thermometer_o[200] sky130_fd_sc_hd__clkbuf_2
Xoutput171 _3263_/X VGND VGND VPWR VPWR output_thermometer_o[135] sky130_fd_sc_hd__clkbuf_2
Xoutput182 _3333_/X VGND VGND VPWR VPWR output_thermometer_o[205] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2150_ _2158_/A _2809_/A VGND VGND VPWR VPWR _3038_/B sky130_fd_sc_hd__and2_1
X_2081_ _2081_/A _2081_/B VGND VGND VPWR VPWR _2784_/B sky130_fd_sc_hd__nor2_4
X_2983_ _2990_/A _2983_/B VGND VGND VPWR VPWR _2983_/X sky130_fd_sc_hd__or2_1
X_1934_ _1934_/A VGND VGND VPWR VPWR _2491_/A sky130_fd_sc_hd__inv_2
X_1865_ _1878_/A _1865_/B VGND VGND VPWR VPWR _1865_/Y sky130_fd_sc_hd__nor2_1
X_1796_ _2961_/A VGND VGND VPWR VPWR _2936_/A sky130_fd_sc_hd__clkbuf_2
X_2417_ _2676_/B _2171_/X _2416_/X VGND VGND VPWR VPWR _2417_/Y sky130_fd_sc_hd__o21ai_1
X_3397_ _3404_/CLK _3397_/D input1/X VGND VGND VPWR VPWR _3398_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2348_ _2347_/X _2022_/A _1988_/A VGND VGND VPWR VPWR _2650_/A sky130_fd_sc_hd__o21a_1
X_2279_ _2279_/A _2286_/B VGND VGND VPWR VPWR _2621_/B sky130_fd_sc_hd__nor2_2
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ _1658_/B VGND VGND VPWR VPWR _2907_/A sky130_fd_sc_hd__inv_2
X_1581_ _2131_/A VGND VGND VPWR VPWR _1581_/X sky130_fd_sc_hd__buf_2
X_3320_ _2174_/Y _2219_/A _3382_/S VGND VGND VPWR VPWR _3320_/X sky130_fd_sc_hd__mux2_2
X_3251_ _3034_/Y _3031_/Y _3380_/S VGND VGND VPWR VPWR _3251_/X sky130_fd_sc_hd__mux2_2
X_3182_ _2786_/Y _2784_/Y _3374_/S VGND VGND VPWR VPWR _3182_/X sky130_fd_sc_hd__mux2_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2202_ _2682_/A VGND VGND VPWR VPWR _2202_/X sky130_fd_sc_hd__clkbuf_2
X_2133_ _2149_/A _2133_/B _2141_/C VGND VGND VPWR VPWR _2803_/A sky130_fd_sc_hd__or3_4
XFILLER_66_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2064_ _2042_/X _2067_/B _2030_/X _2044_/X VGND VGND VPWR VPWR _2070_/B sky130_fd_sc_hd__a31o_1
XFILLER_34_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2966_ _2959_/X _1912_/B _2960_/X _2730_/B _2965_/X VGND VGND VPWR VPWR _2966_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2897_ _2905_/A _2897_/B VGND VGND VPWR VPWR _2897_/Y sky130_fd_sc_hd__nor2_1
X_1917_ _1917_/A _2481_/A _1954_/C VGND VGND VPWR VPWR _1917_/X sky130_fd_sc_hd__or3_1
X_1848_ _2067_/A _2043_/A VGND VGND VPWR VPWR _1849_/A sky130_fd_sc_hd__or2_2
XFILLER_1_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1779_ _1779_/A _1779_/B VGND VGND VPWR VPWR _2697_/B sky130_fd_sc_hd__nor2_2
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2820_ _2820_/A VGND VGND VPWR VPWR _2821_/B sky130_fd_sc_hd__inv_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2751_ _1973_/B _2743_/X _2982_/B _2734_/X _2750_/X VGND VGND VPWR VPWR _2751_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1702_ _2347_/A _1932_/A VGND VGND VPWR VPWR _2124_/B sky130_fd_sc_hd__or2_4
X_2682_ _2682_/A VGND VGND VPWR VPWR _2682_/X sky130_fd_sc_hd__clkbuf_2
X_1633_ _1610_/X _2406_/A _1622_/X _2900_/B VGND VGND VPWR VPWR _1633_/X sky130_fd_sc_hd__o22a_1
X_1564_ _3386_/Q VGND VGND VPWR VPWR _1566_/A sky130_fd_sc_hd__inv_2
X_3303_ _2000_/Y _1996_/Y _3370_/S VGND VGND VPWR VPWR _3303_/X sky130_fd_sc_hd__mux2_2
X_3234_ _2973_/Y _2971_/Y _3383_/S VGND VGND VPWR VPWR _3234_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3165_ _2720_/Y _2718_/Y _3357_/S VGND VGND VPWR VPWR _3165_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2116_ _1755_/X _3024_/B _2114_/B _1802_/X VGND VGND VPWR VPWR _2116_/X sky130_fd_sc_hd__o22a_1
X_3096_ _3107_/A _3096_/B VGND VGND VPWR VPWR _3096_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2047_ _2056_/A _3005_/B VGND VGND VPWR VPWR _2047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2949_ _2956_/A _2949_/B VGND VGND VPWR VPWR _2949_/X sky130_fd_sc_hd__or2_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2803_ _2803_/A _2803_/B VGND VGND VPWR VPWR _2803_/X sky130_fd_sc_hd__or2_1
X_2734_ _2791_/A VGND VGND VPWR VPWR _2734_/X sky130_fd_sc_hd__buf_2
X_2665_ _2606_/X _2894_/B _2664_/X VGND VGND VPWR VPWR _2665_/Y sky130_fd_sc_hd__o21ai_1
X_1616_ _1631_/A _2219_/A VGND VGND VPWR VPWR _2406_/A sky130_fd_sc_hd__nand2_1
X_2596_ _3051_/B _2581_/X _2594_/X _2828_/B _2595_/X VGND VGND VPWR VPWR _2596_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3217_ _2912_/Y _2910_/Y _3346_/S VGND VGND VPWR VPWR _3217_/X sky130_fd_sc_hd__mux2_2
XFILLER_27_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3148_ _2661_/Y _2659_/Y _3340_/S VGND VGND VPWR VPWR _3148_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3079_ _3098_/A VGND VGND VPWR VPWR _3079_/X sky130_fd_sc_hd__buf_2
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2450_ _2514_/B VGND VGND VPWR VPWR _2509_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2381_ _2478_/A VGND VGND VPWR VPWR _2381_/X sky130_fd_sc_hd__buf_2
X_3002_ _2526_/A _2994_/X _2997_/X _2769_/B _3001_/X VGND VGND VPWR VPWR _3002_/Y
+ sky130_fd_sc_hd__o221ai_1
Xinput5 input_binary_i[2] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2717_ _1865_/B _2704_/X _2948_/B _2715_/X _2716_/X VGND VGND VPWR VPWR _2717_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2648_ _3104_/B _2630_/X _1610_/X _2343_/Y _2647_/X VGND VGND VPWR VPWR _2648_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2579_ _2607_/A VGND VGND VPWR VPWR _2766_/A sky130_fd_sc_hd__buf_2
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1950_ _1996_/A _1950_/B VGND VGND VPWR VPWR _1950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1881_ _1917_/A _2467_/A _1893_/C VGND VGND VPWR VPWR _1881_/X sky130_fd_sc_hd__or3_1
X_2502_ _2501_/X _2977_/B _1960_/B _2488_/X VGND VGND VPWR VPWR _2502_/X sky130_fd_sc_hd__o22a_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2433_ _2691_/B _2428_/X _2432_/X VGND VGND VPWR VPWR _2433_/Y sky130_fd_sc_hd__o21ai_1
X_2364_ _2364_/A VGND VGND VPWR VPWR _3111_/B sky130_fd_sc_hd__inv_2
XFILLER_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2295_ _2295_/A _2344_/A VGND VGND VPWR VPWR _2629_/B sky130_fd_sc_hd__nor2_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 _3286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput150 _3379_/X VGND VGND VPWR VPWR output_thermometer_o[251] sky130_fd_sc_hd__clkbuf_2
Xoutput161 _3243_/X VGND VGND VPWR VPWR output_thermometer_o[115] sky130_fd_sc_hd__clkbuf_2
Xoutput183 _3260_/X VGND VGND VPWR VPWR output_thermometer_o[132] sky130_fd_sc_hd__clkbuf_2
Xoutput194 _3232_/X VGND VGND VPWR VPWR output_thermometer_o[104] sky130_fd_sc_hd__clkbuf_2
Xoutput172 _3269_/X VGND VGND VPWR VPWR output_thermometer_o[141] sky130_fd_sc_hd__clkbuf_2
XFILLER_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2080_ _3098_/A VGND VGND VPWR VPWR _2080_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2982_ _2985_/A _2982_/B VGND VGND VPWR VPWR _2982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1933_ _1981_/A _2286_/A VGND VGND VPWR VPWR _1934_/A sky130_fd_sc_hd__or2_2
X_1864_ _1867_/B VGND VGND VPWR VPWR _1865_/B sky130_fd_sc_hd__inv_2
X_1795_ _2993_/A VGND VGND VPWR VPWR _2961_/A sky130_fd_sc_hd__clkbuf_2
X_2416_ _2381_/X _2910_/B _2911_/A _2415_/X VGND VGND VPWR VPWR _2416_/X sky130_fd_sc_hd__o22a_1
X_3396_ _3404_/CLK _3396_/D input1/X VGND VGND VPWR VPWR _3397_/D sky130_fd_sc_hd__dfrtp_1
X_2347_ _2347_/A VGND VGND VPWR VPWR _2347_/X sky130_fd_sc_hd__clkbuf_4
X_2278_ _2279_/A _2317_/B VGND VGND VPWR VPWR _3077_/B sky130_fd_sc_hd__nor2_2
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1580_ _2523_/A VGND VGND VPWR VPWR _2131_/A sky130_fd_sc_hd__buf_2
X_3250_ _3030_/Y _3028_/Y _3381_/S VGND VGND VPWR VPWR _3250_/X sky130_fd_sc_hd__mux2_2
X_3181_ _2783_/Y _2781_/Y _3374_/S VGND VGND VPWR VPWR _3181_/X sky130_fd_sc_hd__mux2_2
X_2201_ _2426_/A VGND VGND VPWR VPWR _2682_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2132_ _2156_/A _2132_/B VGND VGND VPWR VPWR _2802_/B sky130_fd_sc_hd__nor2_2
X_2063_ _3047_/A VGND VGND VPWR VPWR _2109_/A sky130_fd_sc_hd__buf_1
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2965_ _2975_/A _2965_/B VGND VGND VPWR VPWR _2965_/X sky130_fd_sc_hd__or2_1
X_2896_ _1818_/X _2663_/B _2895_/X VGND VGND VPWR VPWR _2896_/Y sky130_fd_sc_hd__o21ai_1
X_1916_ _1964_/A _1916_/B VGND VGND VPWR VPWR _2730_/B sky130_fd_sc_hd__nor2_4
X_1847_ _1847_/A _2057_/A VGND VGND VPWR VPWR _2043_/A sky130_fd_sc_hd__or2_1
X_1778_ _2193_/A VGND VGND VPWR VPWR _1779_/A sky130_fd_sc_hd__buf_4
X_3379_ _2561_/Y _2559_/Y _3381_/S VGND VGND VPWR VPWR _3379_/X sky130_fd_sc_hd__mux2_2
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _2785_/C _2983_/B VGND VGND VPWR VPWR _2750_/X sky130_fd_sc_hd__or2_1
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2681_ _2694_/A _2681_/B VGND VGND VPWR VPWR _2681_/Y sky130_fd_sc_hd__nor2_1
X_1701_ _1808_/B _1833_/A _1744_/A VGND VGND VPWR VPWR _1932_/A sky130_fd_sc_hd__o21ai_2
X_1632_ _1725_/A _1725_/B _1632_/C VGND VGND VPWR VPWR _2900_/B sky130_fd_sc_hd__and3_1
X_3302_ _1990_/Y _1985_/Y _3370_/S VGND VGND VPWR VPWR _3302_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3233_ _2969_/Y _2967_/Y _3365_/S VGND VGND VPWR VPWR _3233_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3164_ _2717_/Y _2714_/Y _3357_/S VGND VGND VPWR VPWR _3164_/X sky130_fd_sc_hd__mux2_1
X_2115_ _2142_/A _2795_/A VGND VGND VPWR VPWR _3024_/B sky130_fd_sc_hd__and2_1
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3095_ _3078_/X _2868_/B _3079_/X _2636_/B _3094_/X VGND VGND VPWR VPWR _3095_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2046_ _2051_/B VGND VGND VPWR VPWR _3005_/B sky130_fd_sc_hd__inv_2
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2948_ _2948_/A _2948_/B VGND VGND VPWR VPWR _2948_/Y sky130_fd_sc_hd__nor2_1
X_2879_ _2887_/A _3107_/B _2879_/C VGND VGND VPWR VPWR _2879_/X sky130_fd_sc_hd__or3_1
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater280 _3351_/S VGND VGND VPWR VPWR _3342_/S sky130_fd_sc_hd__buf_6
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2802_ _2811_/A _2802_/B VGND VGND VPWR VPWR _2802_/Y sky130_fd_sc_hd__nor2_1
X_2733_ _2737_/A _2733_/B VGND VGND VPWR VPWR _2733_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2664_ _2936_/A _3120_/A _2387_/B _2584_/X VGND VGND VPWR VPWR _2664_/X sky130_fd_sc_hd__o22a_1
X_1615_ _2398_/A VGND VGND VPWR VPWR _2219_/A sky130_fd_sc_hd__inv_2
X_2595_ _2705_/A _3054_/B VGND VGND VPWR VPWR _2595_/X sky130_fd_sc_hd__or2_1
X_3216_ _2908_/Y _2905_/Y _3347_/S VGND VGND VPWR VPWR _3216_/X sky130_fd_sc_hd__mux2_1
X_3147_ _2658_/Y _2656_/Y _3357_/S VGND VGND VPWR VPWR _3147_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3078_ _3097_/A VGND VGND VPWR VPWR _3078_/X sky130_fd_sc_hd__buf_2
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2029_ _2029_/A VGND VGND VPWR VPWR _2207_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2380_ _2380_/A _2383_/A VGND VGND VPWR VPWR _2659_/B sky130_fd_sc_hd__nor2_4
X_3001_ _3001_/A _3001_/B VGND VGND VPWR VPWR _3001_/X sky130_fd_sc_hd__or2_1
Xinput6 input_binary_i[3] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2716_ _2724_/A _2949_/B VGND VGND VPWR VPWR _2716_/X sky130_fd_sc_hd__or2_1
X_2647_ _3105_/B _2660_/B VGND VGND VPWR VPWR _2647_/X sky130_fd_sc_hd__or2_1
X_2578_ _2578_/A _2578_/B VGND VGND VPWR VPWR _2607_/A sky130_fd_sc_hd__or2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1903_/A _1880_/B VGND VGND VPWR VPWR _2718_/B sky130_fd_sc_hd__nor2_4
X_2501_ _2523_/A VGND VGND VPWR VPWR _2501_/X sky130_fd_sc_hd__clkbuf_2
X_2432_ _2422_/X _2924_/B _2925_/A _2415_/X VGND VGND VPWR VPWR _2432_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2363_ _2291_/X _2654_/A _2234_/X VGND VGND VPWR VPWR _2881_/B sky130_fd_sc_hd__o21a_1
X_2294_ _2390_/A VGND VGND VPWR VPWR _2294_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _3285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput151 _3290_/X VGND VGND VPWR VPWR output_thermometer_o[162] sky130_fd_sc_hd__clkbuf_2
Xoutput140 _3270_/X VGND VGND VPWR VPWR output_thermometer_o[142] sky130_fd_sc_hd__clkbuf_2
Xoutput173 _3218_/X VGND VGND VPWR VPWR output_thermometer_o[90] sky130_fd_sc_hd__clkbuf_2
Xoutput195 _3264_/X VGND VGND VPWR VPWR output_thermometer_o[136] sky130_fd_sc_hd__clkbuf_2
Xoutput162 _3190_/X VGND VGND VPWR VPWR output_thermometer_o[62] sky130_fd_sc_hd__clkbuf_2
Xoutput184 _3287_/X VGND VGND VPWR VPWR output_thermometer_o[159] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2981_ _2978_/X _1960_/B _2979_/X _2746_/B _2980_/X VGND VGND VPWR VPWR _2981_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1932_ _1932_/A VGND VGND VPWR VPWR _2286_/A sky130_fd_sc_hd__clkinv_4
X_1863_ _1806_/X _2462_/A _2093_/A VGND VGND VPWR VPWR _1867_/B sky130_fd_sc_hd__o21ai_2
X_1794_ _1794_/A VGND VGND VPWR VPWR _1794_/Y sky130_fd_sc_hd__inv_2
X_2415_ _2849_/A VGND VGND VPWR VPWR _2415_/X sky130_fd_sc_hd__clkbuf_2
X_3395_ _3404_/CLK _3395_/D input1/X VGND VGND VPWR VPWR _3396_/D sky130_fd_sc_hd__dfrtp_1
X_2346_ _2173_/X _3104_/B _2345_/X VGND VGND VPWR VPWR _2346_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2277_ _2277_/A VGND VGND VPWR VPWR _2317_/B sky130_fd_sc_hd__buf_2
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2200_ _3054_/B VGND VGND VPWR VPWR _2200_/Y sky130_fd_sc_hd__inv_2
X_3180_ _2778_/Y _2776_/Y _3370_/S VGND VGND VPWR VPWR _3180_/X sky130_fd_sc_hd__mux2_2
X_2131_ _2131_/A VGND VGND VPWR VPWR _2131_/X sky130_fd_sc_hd__buf_2
X_2062_ _2034_/X _3008_/B _2025_/X _2776_/B _2061_/X VGND VGND VPWR VPWR _2062_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2964_ _2967_/A _2964_/B VGND VGND VPWR VPWR _2964_/Y sky130_fd_sc_hd__nor2_1
X_1915_ _2038_/A VGND VGND VPWR VPWR _1964_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2895_ _3054_/A _3120_/A _2341_/X _2388_/A VGND VGND VPWR VPWR _2895_/X sky130_fd_sc_hd__o22a_1
X_1846_ _1818_/X _2938_/B _1842_/X _2707_/B _1845_/X VGND VGND VPWR VPWR _1846_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1777_ _2025_/A VGND VGND VPWR VPWR _1777_/X sky130_fd_sc_hd__buf_2
X_3378_ _2558_/Y _2556_/Y _3380_/S VGND VGND VPWR VPWR _3378_/X sky130_fd_sc_hd__mux2_1
X_2329_ _2401_/A _2329_/B VGND VGND VPWR VPWR _3101_/A sky130_fd_sc_hd__nand2_2
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _2759_/A VGND VGND VPWR VPWR _2694_/A sky130_fd_sc_hd__clkbuf_2
X_1700_ _1759_/B VGND VGND VPWR VPWR _1833_/A sky130_fd_sc_hd__inv_2
X_1631_ _1631_/A _1631_/B VGND VGND VPWR VPWR _1632_/C sky130_fd_sc_hd__nand2_1
X_3301_ _1979_/Y _1973_/Y _3370_/S VGND VGND VPWR VPWR _3301_/X sky130_fd_sc_hd__mux2_2
X_3232_ _2966_/Y _2964_/Y _3383_/S VGND VGND VPWR VPWR _3232_/X sky130_fd_sc_hd__mux2_1
X_3163_ _2713_/Y _2711_/Y _3354_/S VGND VGND VPWR VPWR _3163_/X sky130_fd_sc_hd__mux2_2
X_2114_ _2149_/A _2114_/B _2141_/C VGND VGND VPWR VPWR _2795_/A sky130_fd_sc_hd__or3_4
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3094_ _3099_/A _3094_/B _3094_/C VGND VGND VPWR VPWR _3094_/X sky130_fd_sc_hd__or3_1
X_2045_ _2042_/X _2215_/A _2030_/X _2044_/X VGND VGND VPWR VPWR _2051_/B sky130_fd_sc_hd__a31o_1
X_2947_ _2940_/X _1852_/B _2941_/X _2711_/B _2946_/X VGND VGND VPWR VPWR _2947_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2878_ _2886_/A _2878_/B VGND VGND VPWR VPWR _2878_/Y sky130_fd_sc_hd__nor2_1
X_1829_ _2082_/C VGND VGND VPWR VPWR _3105_/A sky130_fd_sc_hd__buf_2
XFILLER_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater281 _3383_/S VGND VGND VPWR VPWR _3357_/S sky130_fd_sc_hd__buf_6
XFILLER_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2801_ _3029_/B _2799_/X _3028_/B _2791_/X _2800_/X VGND VGND VPWR VPWR _2801_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2732_ _1912_/B _2723_/X _2964_/B _2715_/X _2731_/X VGND VGND VPWR VPWR _2732_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2663_ _2676_/A _2663_/B VGND VGND VPWR VPWR _2663_/Y sky130_fd_sc_hd__nor2_1
X_1614_ _2815_/A VGND VGND VPWR VPWR _2398_/A sky130_fd_sc_hd__clkbuf_2
X_2594_ _2715_/A VGND VGND VPWR VPWR _2594_/X sky130_fd_sc_hd__buf_2
X_3215_ _2904_/Y _2900_/Y _3382_/S VGND VGND VPWR VPWR _3215_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3146_ _2655_/Y _2652_/Y _3340_/S VGND VGND VPWR VPWR _3146_/X sky130_fd_sc_hd__mux2_1
X_3077_ _3083_/A _3077_/B VGND VGND VPWR VPWR _3077_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2028_ _1974_/X _2996_/B _2025_/X _2765_/B _2027_/X VGND VGND VPWR VPWR _2028_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3000_ _3003_/A _3000_/B VGND VGND VPWR VPWR _3000_/Y sky130_fd_sc_hd__nor2_1
Xinput7 input_binary_i[4] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2715_ _2715_/A VGND VGND VPWR VPWR _2715_/X sky130_fd_sc_hd__clkbuf_2
X_2646_ _2792_/B VGND VGND VPWR VPWR _2660_/B sky130_fd_sc_hd__buf_1
X_2577_ _2577_/A _2577_/B VGND VGND VPWR VPWR _3354_/S sky130_fd_sc_hd__nor2_8
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3129_ _2591_/Y _2588_/Y _3330_/S VGND VGND VPWR VPWR _3129_/X sky130_fd_sc_hd__mux2_2
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2500_ _2980_/B VGND VGND VPWR VPWR _2500_/Y sky130_fd_sc_hd__inv_2
X_2431_ _2431_/A VGND VGND VPWR VPWR _2431_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2362_ _2380_/A _2364_/A VGND VGND VPWR VPWR _2652_/B sky130_fd_sc_hd__nor2_2
X_2293_ _2295_/A _2317_/B VGND VGND VPWR VPWR _3087_/B sky130_fd_sc_hd__nor2_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_12 _3342_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput152 _3138_/X VGND VGND VPWR VPWR output_thermometer_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput130 _3267_/X VGND VGND VPWR VPWR output_thermometer_o[139] sky130_fd_sc_hd__clkbuf_2
Xoutput141 _3327_/X VGND VGND VPWR VPWR output_thermometer_o[199] sky130_fd_sc_hd__clkbuf_2
X_2629_ _2636_/A _2629_/B VGND VGND VPWR VPWR _2629_/Y sky130_fd_sc_hd__nor2_1
Xoutput174 _3130_/X VGND VGND VPWR VPWR output_thermometer_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput163 _3297_/X VGND VGND VPWR VPWR output_thermometer_o[169] sky130_fd_sc_hd__clkbuf_2
Xoutput185 _3160_/X VGND VGND VPWR VPWR output_thermometer_o[32] sky130_fd_sc_hd__clkbuf_2
Xoutput196 _3161_/X VGND VGND VPWR VPWR output_thermometer_o[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2980_ _2990_/A _2980_/B VGND VGND VPWR VPWR _2980_/X sky130_fd_sc_hd__or2_1
X_1931_ _2157_/A VGND VGND VPWR VPWR _1931_/X sky130_fd_sc_hd__buf_2
X_1862_ _2221_/B VGND VGND VPWR VPWR _2462_/A sky130_fd_sc_hd__inv_2
Xinput10 input_binary_i[7] VGND VGND VPWR VPWR _3389_/D sky130_fd_sc_hd__clkbuf_1
X_1793_ _1988_/A _1792_/Y _2841_/A VGND VGND VPWR VPWR _1794_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2414_ _2435_/A VGND VGND VPWR VPWR _2849_/A sky130_fd_sc_hd__buf_2
X_3394_ _3404_/CLK _3394_/D input1/X VGND VGND VPWR VPWR _3395_/D sky130_fd_sc_hd__dfrtp_1
X_2345_ _2341_/X _2343_/Y _2294_/X _2645_/B VGND VGND VPWR VPWR _2345_/X sky130_fd_sc_hd__o22a_1
X_2276_ _2184_/X _3081_/B _2185_/X VGND VGND VPWR VPWR _2853_/B sky130_fd_sc_hd__o21a_1
XFILLER_52_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2130_ _2155_/A _3033_/B VGND VGND VPWR VPWR _2130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2061_ _2534_/A _2061_/B VGND VGND VPWR VPWR _2061_/X sky130_fd_sc_hd__or2_1
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2963_ _2959_/X _1899_/B _2960_/X _2726_/B _2962_/X VGND VGND VPWR VPWR _2963_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1914_ _1890_/X _1909_/A _1900_/X VGND VGND VPWR VPWR _2964_/B sky130_fd_sc_hd__a21oi_4
X_2894_ _2905_/A _2894_/B VGND VGND VPWR VPWR _2894_/Y sky130_fd_sc_hd__nor2_1
X_1845_ _1858_/A _2452_/A _1893_/C VGND VGND VPWR VPWR _1845_/X sky130_fd_sc_hd__or3_2
X_1776_ _2523_/A VGND VGND VPWR VPWR _2025_/A sky130_fd_sc_hd__clkbuf_2
X_3377_ _2555_/Y _2553_/Y _3381_/S VGND VGND VPWR VPWR _3377_/X sky130_fd_sc_hd__mux2_2
X_2328_ _2727_/A VGND VGND VPWR VPWR _2328_/X sky130_fd_sc_hd__buf_2
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2259_ _2841_/A VGND VGND VPWR VPWR _3110_/A sky130_fd_sc_hd__buf_2
XFILLER_13_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _2044_/A VGND VGND VPWR VPWR _1631_/B sky130_fd_sc_hd__clkbuf_4
X_3300_ _1967_/Y _1960_/Y _3365_/S VGND VGND VPWR VPWR _3300_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3231_ _2963_/Y _2958_/Y _3365_/S VGND VGND VPWR VPWR _3231_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3162_ _2710_/Y _2707_/Y _3354_/S VGND VGND VPWR VPWR _3162_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2113_ _2113_/A VGND VGND VPWR VPWR _2149_/A sky130_fd_sc_hd__buf_1
XFILLER_66_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3093_ _3107_/A _3093_/B VGND VGND VPWR VPWR _3093_/Y sky130_fd_sc_hd__nor2_1
X_2044_ _2044_/A VGND VGND VPWR VPWR _2044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2946_ _2956_/A _2946_/B VGND VGND VPWR VPWR _2946_/X sky130_fd_sc_hd__or2_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2877_ _2851_/A _2339_/Y _2340_/A _2820_/A _2849_/Y VGND VGND VPWR VPWR _2877_/X
+ sky130_fd_sc_hd__a221o_1
X_1828_ _2009_/C VGND VGND VPWR VPWR _2082_/C sky130_fd_sc_hd__clkbuf_2
X_1759_ _1759_/A _1759_/B VGND VGND VPWR VPWR _1884_/B sky130_fd_sc_hd__or2_1
XFILLER_38_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater271 _3342_/S VGND VGND VPWR VPWR _3346_/S sky130_fd_sc_hd__buf_8
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater282 _3354_/S VGND VGND VPWR VPWR _3383_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2800_ _2800_/A _2803_/B VGND VGND VPWR VPWR _2800_/X sky130_fd_sc_hd__or2_1
X_2731_ _2744_/A _2965_/B VGND VGND VPWR VPWR _2731_/X sky130_fd_sc_hd__or2_1
XFILLER_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2662_ _2662_/A VGND VGND VPWR VPWR _2676_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1613_ _1827_/B VGND VGND VPWR VPWR _2815_/A sky130_fd_sc_hd__clkbuf_2
X_2593_ _2610_/A _2593_/B VGND VGND VPWR VPWR _2593_/Y sky130_fd_sc_hd__nor2_1
X_3214_ _2899_/Y _2897_/Y _3342_/S VGND VGND VPWR VPWR _3214_/X sky130_fd_sc_hd__mux2_2
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3145_ _2651_/Y _2649_/Y _3357_/S VGND VGND VPWR VPWR _3145_/X sky130_fd_sc_hd__mux2_1
X_3076_ _3105_/A _2618_/A _2097_/X _2271_/Y _3075_/X VGND VGND VPWR VPWR _3076_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2027_ _2522_/A _2061_/B VGND VGND VPWR VPWR _2027_/X sky130_fd_sc_hd__or2_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2929_ _2929_/A _2939_/A VGND VGND VPWR VPWR _2929_/X sky130_fd_sc_hd__or2_1
XFILLER_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 input_binary_i[5] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2714_ _2718_/A _2714_/B VGND VGND VPWR VPWR _2714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2645_ _2931_/A _2645_/B VGND VGND VPWR VPWR _2645_/Y sky130_fd_sc_hd__nor2_1
X_2576_ _2574_/Y _2575_/Y _2574_/Y _2575_/Y VGND VGND VPWR VPWR _3394_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3128_ _2585_/Y _1725_/B _3382_/S VGND VGND VPWR VPWR _3128_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3059_ _3052_/X _2831_/B _3053_/X _2597_/B _3058_/X VGND VGND VPWR VPWR _3059_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2430_ _2688_/B _2428_/X _2429_/X VGND VGND VPWR VPWR _2430_/Y sky130_fd_sc_hd__o21ai_1
X_2361_ _1639_/X _2036_/A _1648_/A VGND VGND VPWR VPWR _2364_/A sky130_fd_sc_hd__o21ai_2
X_2292_ _2291_/X _3088_/B _2185_/X VGND VGND VPWR VPWR _2861_/B sky130_fd_sc_hd__o21a_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput131 _3376_/X VGND VGND VPWR VPWR output_thermometer_o[248] sky130_fd_sc_hd__clkbuf_2
X_2628_ _3083_/B _2602_/X _2626_/X _2856_/B _2627_/X VGND VGND VPWR VPWR _2628_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput120 _3374_/X VGND VGND VPWR VPWR output_thermometer_o[246] sky130_fd_sc_hd__clkbuf_2
Xoutput142 _3368_/X VGND VGND VPWR VPWR output_thermometer_o[240] sky130_fd_sc_hd__clkbuf_2
X_2559_ _2565_/A _2803_/A VGND VGND VPWR VPWR _2559_/Y sky130_fd_sc_hd__nor2_1
Xoutput153 _3134_/X VGND VGND VPWR VPWR output_thermometer_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput175 _3341_/X VGND VGND VPWR VPWR output_thermometer_o[213] sky130_fd_sc_hd__clkbuf_2
Xoutput164 _3133_/X VGND VGND VPWR VPWR output_thermometer_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput186 _3361_/X VGND VGND VPWR VPWR output_thermometer_o[233] sky130_fd_sc_hd__clkbuf_2
Xoutput197 _3302_/X VGND VGND VPWR VPWR output_thermometer_o[174] sky130_fd_sc_hd__clkbuf_2
XFILLER_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1930_ _1913_/X _2967_/B _1902_/X _2733_/B _1929_/X VGND VGND VPWR VPWR _1930_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1861_ _1907_/A _2057_/A VGND VGND VPWR VPWR _2221_/B sky130_fd_sc_hd__or2_4
Xinput11 input_binary_i[8] VGND VGND VPWR VPWR _3390_/D sky130_fd_sc_hd__clkbuf_1
X_1792_ _1792_/A VGND VGND VPWR VPWR _1792_/Y sky130_fd_sc_hd__inv_2
X_2413_ _2413_/A VGND VGND VPWR VPWR _2413_/Y sky130_fd_sc_hd__inv_2
X_3393_ _3404_/CLK input4/X VGND VGND VPWR VPWR _3393_/Q sky130_fd_sc_hd__dfxtp_2
X_2344_ _2344_/A VGND VGND VPWR VPWR _2645_/B sky130_fd_sc_hd__inv_2
X_2275_ _2290_/A _3081_/B VGND VGND VPWR VPWR _2275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2060_ _2081_/A _2060_/B VGND VGND VPWR VPWR _2776_/B sky130_fd_sc_hd__nor2_4
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2962_ _2975_/A _2962_/B VGND VGND VPWR VPWR _2962_/X sky130_fd_sc_hd__or2_1
X_1913_ _2087_/A VGND VGND VPWR VPWR _1913_/X sky130_fd_sc_hd__buf_2
X_2893_ _2882_/X _2659_/B _2331_/X _3118_/B _2892_/X VGND VGND VPWR VPWR _2893_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1844_ _2082_/C VGND VGND VPWR VPWR _1893_/C sky130_fd_sc_hd__buf_1
X_1775_ _1786_/A _2440_/A VGND VGND VPWR VPWR _1775_/Y sky130_fd_sc_hd__nor2_1
X_3376_ _2551_/Y _2548_/Y _3381_/S VGND VGND VPWR VPWR _3376_/X sky130_fd_sc_hd__mux2_1
X_2327_ _2617_/B VGND VGND VPWR VPWR _2327_/Y sky130_fd_sc_hd__inv_2
X_2258_ _3044_/A _2262_/A VGND VGND VPWR VPWR _2258_/Y sky130_fd_sc_hd__nor2_1
X_2189_ _3390_/Q _2189_/B VGND VGND VPWR VPWR _2277_/A sky130_fd_sc_hd__or2_2
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _2957_/Y _2955_/Y _3383_/S VGND VGND VPWR VPWR _3230_/X sky130_fd_sc_hd__mux2_2
X_3161_ _2706_/Y _2703_/Y _3354_/S VGND VGND VPWR VPWR _3161_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2112_ _2234_/A VGND VGND VPWR VPWR _2142_/A sky130_fd_sc_hd__clkbuf_2
X_3092_ _3078_/X _2864_/B _3079_/X _2633_/B _3091_/X VGND VGND VPWR VPWR _3092_/Y
+ sky130_fd_sc_hd__o221ai_2
X_2043_ _2043_/A VGND VGND VPWR VPWR _2215_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2945_ _2948_/A _2945_/B VGND VGND VPWR VPWR _2945_/Y sky130_fd_sc_hd__nor2_1
X_2876_ _2324_/X _3101_/A _2875_/X VGND VGND VPWR VPWR _2876_/Y sky130_fd_sc_hd__o21ai_1
X_1827_ _2168_/A _1827_/B VGND VGND VPWR VPWR _2009_/C sky130_fd_sc_hd__or2_1
X_1758_ _1735_/X _2691_/B _1757_/X VGND VGND VPWR VPWR _1758_/Y sky130_fd_sc_hd__o21ai_1
X_1689_ _2089_/A _1689_/B VGND VGND VPWR VPWR _2676_/B sky130_fd_sc_hd__nor2_4
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3359_ _2480_/Y _2477_/Y _3383_/S VGND VGND VPWR VPWR _3359_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater272 _3382_/S VGND VGND VPWR VPWR _3381_/S sky130_fd_sc_hd__buf_8
Xrepeater283 _3354_/S VGND VGND VPWR VPWR _3351_/S sky130_fd_sc_hd__buf_8
XFILLER_53_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2730_ _2737_/A _2730_/B VGND VGND VPWR VPWR _2730_/Y sky130_fd_sc_hd__nor2_1
X_2661_ _3117_/B _2653_/X _2171_/A _2891_/B _2660_/X VGND VGND VPWR VPWR _2661_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1612_ _2101_/A _1588_/Y _1642_/A _2161_/A VGND VGND VPWR VPWR _1827_/B sky130_fd_sc_hd__a31o_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2592_ _2662_/A VGND VGND VPWR VPWR _2610_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3213_ _2896_/Y _2894_/Y _3382_/S VGND VGND VPWR VPWR _3213_/X sky130_fd_sc_hd__mux2_1
X_3144_ _2648_/Y _2645_/Y _3354_/S VGND VGND VPWR VPWR _3144_/X sky130_fd_sc_hd__mux2_1
X_3075_ _2301_/C _2269_/A _2131_/A VGND VGND VPWR VPWR _3075_/X sky130_fd_sc_hd__a21o_1
X_2026_ _2026_/A _2026_/B VGND VGND VPWR VPWR _2765_/B sky130_fd_sc_hd__nor2_2
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2928_ _2948_/A _2928_/B VGND VGND VPWR VPWR _2928_/Y sky130_fd_sc_hd__nor2_1
X_2859_ _3084_/B _2932_/B VGND VGND VPWR VPWR _2859_/X sky130_fd_sc_hd__or2_1
XFILLER_49_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 input_binary_i[6] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2713_ _1852_/B _2704_/X _2945_/B _2673_/X _2712_/X VGND VGND VPWR VPWR _2713_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2644_ _2324_/X _2335_/Y _2643_/X VGND VGND VPWR VPWR _2644_/Y sky130_fd_sc_hd__o21ai_1
X_2575_ _3396_/D _3395_/D _3396_/D _3395_/D VGND VGND VPWR VPWR _2575_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3127_ VGND VGND VPWR VPWR _3127_/HI _3383_/A1 sky130_fd_sc_hd__conb_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3058_ _3058_/A _3058_/B _3094_/C VGND VGND VPWR VPWR _3058_/X sky130_fd_sc_hd__or3_1
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2009_ _2103_/A _2009_/B _2009_/C VGND VGND VPWR VPWR _2090_/B sky130_fd_sc_hd__or3_1
XFILLER_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ _3112_/B VGND VGND VPWR VPWR _2360_/Y sky130_fd_sc_hd__inv_2
X_2291_ _2291_/A VGND VGND VPWR VPWR _2291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput110 _3132_/X VGND VGND VPWR VPWR output_thermometer_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput121 _3281_/X VGND VGND VPWR VPWR output_thermometer_o[153] sky130_fd_sc_hd__clkbuf_2
Xoutput143 _3231_/X VGND VGND VPWR VPWR output_thermometer_o[103] sky130_fd_sc_hd__clkbuf_2
X_2627_ _3084_/B _2641_/B VGND VGND VPWR VPWR _2627_/X sky130_fd_sc_hd__or2_1
Xoutput132 _3318_/X VGND VGND VPWR VPWR output_thermometer_o[190] sky130_fd_sc_hd__clkbuf_2
X_2558_ _2315_/X _3028_/B _2557_/X VGND VGND VPWR VPWR _2558_/Y sky130_fd_sc_hd__o21ai_1
Xoutput165 _3268_/X VGND VGND VPWR VPWR output_thermometer_o[140] sky130_fd_sc_hd__clkbuf_2
Xoutput176 _3221_/X VGND VGND VPWR VPWR output_thermometer_o[93] sky130_fd_sc_hd__clkbuf_2
Xoutput154 _3276_/X VGND VGND VPWR VPWR output_thermometer_o[148] sky130_fd_sc_hd__clkbuf_2
Xoutput198 _3337_/X VGND VGND VPWR VPWR output_thermometer_o[209] sky130_fd_sc_hd__clkbuf_2
Xoutput187 _3336_/X VGND VGND VPWR VPWR output_thermometer_o[208] sky130_fd_sc_hd__clkbuf_2
X_2489_ _2478_/X _2967_/B _1925_/B _2488_/X VGND VGND VPWR VPWR _2489_/X sky130_fd_sc_hd__o22a_1
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ _1860_/A VGND VGND VPWR VPWR _1907_/A sky130_fd_sc_hd__buf_1
X_1791_ _3391_/Q _1791_/B VGND VGND VPWR VPWR _1792_/A sky130_fd_sc_hd__or2_2
Xinput12 input_binary_i[9] VGND VGND VPWR VPWR _3391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2412_ _2315_/X _2905_/B _2411_/X VGND VGND VPWR VPWR _2412_/Y sky130_fd_sc_hd__o21ai_1
X_3392_ _3408_/CLK input3/X VGND VGND VPWR VPWR _3392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2343_ _2343_/A VGND VGND VPWR VPWR _2343_/Y sky130_fd_sc_hd__inv_2
X_2274_ _2279_/A _2289_/B VGND VGND VPWR VPWR _3081_/B sky130_fd_sc_hd__nor2_2
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1989_ _2082_/A _2509_/A _2071_/C VGND VGND VPWR VPWR _1989_/X sky130_fd_sc_hd__or3_1
XFILLER_57_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2961_ _2961_/A VGND VGND VPWR VPWR _2975_/A sky130_fd_sc_hd__buf_1
X_1912_ _1938_/A _1912_/B VGND VGND VPWR VPWR _1912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2892_ _2898_/A _3117_/B _3049_/C VGND VGND VPWR VPWR _2892_/X sky130_fd_sc_hd__or3_1
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1843_ _3044_/A _1843_/B VGND VGND VPWR VPWR _2707_/B sky130_fd_sc_hd__nor2_2
X_1774_ _1779_/B VGND VGND VPWR VPWR _2440_/A sky130_fd_sc_hd__inv_2
X_3375_ _2547_/Y _3019_/B _3381_/S VGND VGND VPWR VPWR _3375_/X sky130_fd_sc_hd__mux2_1
X_2326_ _2326_/A VGND VGND VPWR VPWR _2617_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2257_ _2257_/A _2329_/B VGND VGND VPWR VPWR _2262_/A sky130_fd_sc_hd__or2_2
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2188_ _2549_/A VGND VGND VPWR VPWR _2188_/X sky130_fd_sc_hd__buf_2
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3160_ _2701_/Y _1799_/A _3382_/S VGND VGND VPWR VPWR _3160_/X sky130_fd_sc_hd__mux2_1
X_2111_ _2156_/A _2111_/B VGND VGND VPWR VPWR _2794_/B sky130_fd_sc_hd__nor2_2
X_3091_ _3108_/A _3091_/B VGND VGND VPWR VPWR _3091_/X sky130_fd_sc_hd__or2_1
X_2042_ _2042_/A VGND VGND VPWR VPWR _2042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2944_ _2940_/X _1838_/B _2941_/X _2707_/B _2943_/X VGND VGND VPWR VPWR _2944_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2875_ _2328_/X _2327_/Y _2331_/X _2322_/A VGND VGND VPWR VPWR _2875_/X sky130_fd_sc_hd__o22a_1
X_1826_ _1928_/A VGND VGND VPWR VPWR _1858_/A sky130_fd_sc_hd__clkbuf_2
X_1757_ _1708_/X _2431_/A _1755_/X _2924_/B VGND VGND VPWR VPWR _1757_/X sky130_fd_sc_hd__o22a_1
X_1688_ _2038_/A VGND VGND VPWR VPWR _2089_/A sky130_fd_sc_hd__buf_4
X_3358_ _2474_/Y _2472_/Y _3383_/S VGND VGND VPWR VPWR _3358_/X sky130_fd_sc_hd__mux2_4
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2309_ _2310_/A _2317_/B VGND VGND VPWR VPWR _3093_/B sky130_fd_sc_hd__nor2_2
X_3289_ _1831_/Y _1816_/Y _3351_/S VGND VGND VPWR VPWR _3289_/X sky130_fd_sc_hd__mux2_2
Xrepeater273 _3374_/S VGND VGND VPWR VPWR _3370_/S sky130_fd_sc_hd__buf_8
Xrepeater284 _3354_/S VGND VGND VPWR VPWR _3365_/S sky130_fd_sc_hd__buf_8
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2660_ _2660_/A _2660_/B VGND VGND VPWR VPWR _2660_/X sky130_fd_sc_hd__or2_1
X_1611_ _3391_/Q _3390_/Q VGND VGND VPWR VPWR _2161_/A sky130_fd_sc_hd__nand2_2
X_2591_ _3048_/B _2581_/X _2256_/X _2823_/B _2590_/X VGND VGND VPWR VPWR _2591_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3212_ _2893_/Y _2891_/Y _3340_/S VGND VGND VPWR VPWR _3212_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3143_ _2644_/Y _2617_/B _3351_/S VGND VGND VPWR VPWR _3143_/X sky130_fd_sc_hd__mux2_2
X_3074_ _3083_/A _3074_/B VGND VGND VPWR VPWR _3074_/Y sky130_fd_sc_hd__nor2_1
X_2025_ _2025_/A VGND VGND VPWR VPWR _2025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2927_ _2970_/A VGND VGND VPWR VPWR _2948_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2858_ _3022_/B VGND VGND VPWR VPWR _2932_/B sky130_fd_sc_hd__clkbuf_2
X_2789_ _2086_/B _2761_/X _3018_/B _2773_/X _2788_/X VGND VGND VPWR VPWR _2789_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1809_ _3385_/Q _1809_/B _1832_/A VGND VGND VPWR VPWR _2012_/A sky130_fd_sc_hd__or3_4
XFILLER_65_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2712_ _2724_/A _2946_/B VGND VGND VPWR VPWR _2712_/X sky130_fd_sc_hd__or2_1
X_2643_ _2341_/X _3101_/A _2393_/X _2322_/A VGND VGND VPWR VPWR _2643_/X sky130_fd_sc_hd__o22a_1
X_2574_ _3399_/D VGND VGND VPWR VPWR _2574_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3126_ _3126_/A _3126_/B VGND VGND VPWR VPWR _3126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3057_ _3057_/A VGND VGND VPWR VPWR _3094_/C sky130_fd_sc_hd__buf_1
X_2008_ _2347_/A VGND VGND VPWR VPWR _2103_/A sky130_fd_sc_hd__buf_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2290_ _2290_/A _3088_/B VGND VGND VPWR VPWR _2290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2626_ _2715_/A VGND VGND VPWR VPWR _2626_/X sky130_fd_sc_hd__clkbuf_2
Xoutput100 _3191_/X VGND VGND VPWR VPWR output_thermometer_o[63] sky130_fd_sc_hd__clkbuf_2
Xoutput133 _3237_/X VGND VGND VPWR VPWR output_thermometer_o[109] sky130_fd_sc_hd__clkbuf_2
Xoutput111 _3347_/X VGND VGND VPWR VPWR output_thermometer_o[219] sky130_fd_sc_hd__clkbuf_2
Xoutput122 _3282_/X VGND VGND VPWR VPWR output_thermometer_o[154] sky130_fd_sc_hd__clkbuf_2
X_2557_ _2798_/B _2390_/X _3029_/B _2549_/X VGND VGND VPWR VPWR _2557_/X sky130_fd_sc_hd__o22a_1
Xoutput155 _3238_/X VGND VGND VPWR VPWR output_thermometer_o[110] sky130_fd_sc_hd__clkbuf_2
Xoutput177 _3301_/X VGND VGND VPWR VPWR output_thermometer_o[173] sky130_fd_sc_hd__clkbuf_2
Xoutput144 _3266_/X VGND VGND VPWR VPWR output_thermometer_o[138] sky130_fd_sc_hd__clkbuf_2
Xoutput166 _3177_/X VGND VGND VPWR VPWR output_thermometer_o[49] sky130_fd_sc_hd__clkbuf_2
Xoutput199 _3334_/X VGND VGND VPWR VPWR output_thermometer_o[206] sky130_fd_sc_hd__clkbuf_2
X_2488_ _2531_/A VGND VGND VPWR VPWR _2488_/X sky130_fd_sc_hd__clkbuf_2
Xoutput188 _3144_/X VGND VGND VPWR VPWR output_thermometer_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3109_ _3097_/X _2878_/B _3098_/X _2649_/B _3108_/X VGND VGND VPWR VPWR _3109_/Y
+ sky130_fd_sc_hd__o221ai_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1790_ _2092_/C VGND VGND VPWR VPWR _1988_/A sky130_fd_sc_hd__buf_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2411_ _2907_/A _2188_/X _2672_/B _2171_/A VGND VGND VPWR VPWR _2411_/X sky130_fd_sc_hd__o22a_1
X_3391_ _3408_/CLK _3391_/D VGND VGND VPWR VPWR _3391_/Q sky130_fd_sc_hd__dfxtp_2
X_2342_ _2014_/X _1627_/A _2189_/B _2193_/A VGND VGND VPWR VPWR _2343_/A sky130_fd_sc_hd__a31o_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2273_ _2173_/X _3074_/B _1797_/X _2271_/Y _2272_/X VGND VGND VPWR VPWR _2273_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ _1988_/A VGND VGND VPWR VPWR _2082_/A sky130_fd_sc_hd__clkbuf_2
X_2609_ _2606_/X _2839_/B _2608_/X VGND VGND VPWR VPWR _2609_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2960_ _2960_/A VGND VGND VPWR VPWR _2960_/X sky130_fd_sc_hd__buf_2
X_2891_ _2905_/A _2891_/B VGND VGND VPWR VPWR _2891_/Y sky130_fd_sc_hd__nor2_1
X_1911_ _1916_/B VGND VGND VPWR VPWR _1912_/B sky130_fd_sc_hd__inv_2
XFILLER_63_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1842_ _2025_/A VGND VGND VPWR VPWR _1842_/X sky130_fd_sc_hd__buf_2
X_1773_ _2165_/B _1773_/B VGND VGND VPWR VPWR _1779_/B sky130_fd_sc_hd__or2_2
X_3374_ _2543_/Y _3016_/B _3374_/S VGND VGND VPWR VPWR _3374_/X sky130_fd_sc_hd__mux2_2
X_2325_ _2333_/A _2329_/B VGND VGND VPWR VPWR _2326_/A sky130_fd_sc_hd__or2_1
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2256_ _2715_/A VGND VGND VPWR VPWR _2256_/X sky130_fd_sc_hd__buf_2
XFILLER_57_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2187_ _2435_/A VGND VGND VPWR VPWR _2549_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2110_ _2242_/A VGND VGND VPWR VPWR _2156_/A sky130_fd_sc_hd__clkbuf_4
X_3090_ _3090_/A VGND VGND VPWR VPWR _3090_/Y sky130_fd_sc_hd__inv_2
X_2041_ _2034_/X _3000_/B _2025_/X _2769_/B _2040_/X VGND VGND VPWR VPWR _2041_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2943_ _2956_/A _2943_/B VGND VGND VPWR VPWR _2943_/X sky130_fd_sc_hd__or2_1
X_2874_ _2857_/X _3096_/B _2872_/X _2640_/B _2873_/X VGND VGND VPWR VPWR _2874_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1825_ _2009_/B VGND VGND VPWR VPWR _1928_/A sky130_fd_sc_hd__buf_2
X_1756_ _1769_/A _1769_/B _1756_/C VGND VGND VPWR VPWR _2924_/B sky130_fd_sc_hd__and3_1
X_1687_ _2333_/A VGND VGND VPWR VPWR _2038_/A sky130_fd_sc_hd__clkbuf_2
X_3357_ _2470_/Y _2468_/Y _3357_/S VGND VGND VPWR VPWR _3357_/X sky130_fd_sc_hd__mux2_2
X_2308_ _2291_/X _3094_/B _2837_/A VGND VGND VPWR VPWR _2868_/B sky130_fd_sc_hd__o21a_1
X_3288_ _1803_/Y _1786_/Y _3381_/S VGND VGND VPWR VPWR _3288_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater274 _3382_/S VGND VGND VPWR VPWR _3374_/S sky130_fd_sc_hd__buf_8
XFILLER_38_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2239_ _2239_/A _2243_/B VGND VGND VPWR VPWR _2240_/B sky130_fd_sc_hd__nor2_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1610_ _3099_/C VGND VGND VPWR VPWR _1610_/X sky130_fd_sc_hd__buf_2
X_2590_ _3049_/B _2618_/B VGND VGND VPWR VPWR _2590_/X sky130_fd_sc_hd__or2_1
X_3211_ _2888_/Y _2886_/Y _3340_/S VGND VGND VPWR VPWR _3211_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3142_ _2642_/Y _2640_/Y _3340_/S VGND VGND VPWR VPWR _3142_/X sky130_fd_sc_hd__mux2_2
X_3073_ _1777_/X _2258_/Y _3032_/X _2848_/B _3072_/X VGND VGND VPWR VPWR _3073_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2024_ _1992_/X _2019_/X _2020_/X _2522_/A _2023_/X VGND VGND VPWR VPWR _2996_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2926_ _1756_/C _2920_/X _2921_/X _2691_/B _2925_/X VGND VGND VPWR VPWR _2926_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_50_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2857_ _2857_/A VGND VGND VPWR VPWR _2857_/X sky130_fd_sc_hd__buf_2
X_1808_ _3387_/Q _1808_/B VGND VGND VPWR VPWR _1832_/A sky130_fd_sc_hd__or2_1
X_2788_ _2788_/A _2788_/B VGND VGND VPWR VPWR _2788_/X sky130_fd_sc_hd__or2_1
X_1739_ _2185_/A _1740_/C VGND VGND VPWR VPWR _2425_/A sky130_fd_sc_hd__or2_2
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2711_ _2718_/A _2711_/B VGND VGND VPWR VPWR _2711_/Y sky130_fd_sc_hd__nor2_1
X_2642_ _3096_/B _2630_/X _2626_/X _2871_/B _2641_/X VGND VGND VPWR VPWR _2642_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2573_ _2577_/B _2571_/X _2577_/A _2161_/Y VGND VGND VPWR VPWR _2573_/X sky130_fd_sc_hd__a22o_1
X_3125_ _1660_/X _2897_/B _2131_/A _2666_/B _3124_/X VGND VGND VPWR VPWR _3125_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3056_ _3064_/A _3056_/B VGND VGND VPWR VPWR _3056_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2007_ _2026_/A _2007_/B VGND VGND VPWR VPWR _2760_/B sky130_fd_sc_hd__nor2_4
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2909_ _2970_/A VGND VGND VPWR VPWR _2924_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput101 _3137_/X VGND VGND VPWR VPWR output_thermometer_o[9] sky130_fd_sc_hd__clkbuf_2
X_2625_ _2636_/A _2625_/B VGND VGND VPWR VPWR _2625_/Y sky130_fd_sc_hd__nor2_1
Xoutput112 _3128_/X VGND VGND VPWR VPWR output_thermometer_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput123 _3283_/X VGND VGND VPWR VPWR output_thermometer_o[155] sky130_fd_sc_hd__clkbuf_2
Xoutput134 _3209_/X VGND VGND VPWR VPWR output_thermometer_o[81] sky130_fd_sc_hd__clkbuf_2
X_2556_ _2565_/A _2800_/A VGND VGND VPWR VPWR _2556_/Y sky130_fd_sc_hd__nor2_1
Xoutput167 _3277_/X VGND VGND VPWR VPWR output_thermometer_o[149] sky130_fd_sc_hd__clkbuf_2
Xoutput145 _3225_/X VGND VGND VPWR VPWR output_thermometer_o[97] sky130_fd_sc_hd__clkbuf_2
Xoutput156 _3226_/X VGND VGND VPWR VPWR output_thermometer_o[98] sky130_fd_sc_hd__clkbuf_2
Xoutput189 _3291_/X VGND VGND VPWR VPWR output_thermometer_o[163] sky130_fd_sc_hd__clkbuf_2
X_2487_ _2968_/B VGND VGND VPWR VPWR _2487_/Y sky130_fd_sc_hd__inv_2
Xoutput178 _3183_/X VGND VGND VPWR VPWR output_thermometer_o[55] sky130_fd_sc_hd__clkbuf_2
X_3108_ _3108_/A _3108_/B VGND VGND VPWR VPWR _3108_/X sky130_fd_sc_hd__or2_1
X_3039_ _3042_/A _3039_/B VGND VGND VPWR VPWR _3039_/X sky130_fd_sc_hd__or2_1
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2410_ _2410_/A _2674_/A VGND VGND VPWR VPWR _2410_/Y sky130_fd_sc_hd__nor2_1
X_3390_ _3408_/CLK _3390_/D VGND VGND VPWR VPWR _3390_/Q sky130_fd_sc_hd__dfxtp_2
X_2341_ _2961_/A VGND VGND VPWR VPWR _2341_/X sky130_fd_sc_hd__buf_2
X_2272_ _2301_/C _3074_/B _2682_/A VGND VGND VPWR VPWR _2272_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1987_ _2026_/A _1987_/B VGND VGND VPWR VPWR _2752_/B sky130_fd_sc_hd__nor2_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2608_ _3064_/B _2607_/X _2229_/B _2584_/X VGND VGND VPWR VPWR _2608_/X sky130_fd_sc_hd__o22a_1
X_2539_ _2523_/X _3011_/B _3012_/B _2531_/X VGND VGND VPWR VPWR _2539_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2890_ _2970_/A VGND VGND VPWR VPWR _2905_/A sky130_fd_sc_hd__buf_2
X_1910_ _1871_/X _2481_/A _1875_/X VGND VGND VPWR VPWR _1916_/B sky130_fd_sc_hd__o21ai_2
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1841_ _1820_/X _1835_/A _1840_/X VGND VGND VPWR VPWR _2938_/B sky130_fd_sc_hd__a21oi_4
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1772_ _3390_/Q VGND VGND VPWR VPWR _2165_/B sky130_fd_sc_hd__clkbuf_2
X_3373_ _2540_/Y _2538_/Y _3381_/S VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__mux2_4
X_2324_ _3054_/A VGND VGND VPWR VPWR _2324_/X sky130_fd_sc_hd__buf_2
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2255_ _2390_/A VGND VGND VPWR VPWR _2715_/A sky130_fd_sc_hd__clkbuf_2
X_2186_ _2184_/X _3049_/B _2185_/X VGND VGND VPWR VPWR _2823_/B sky130_fd_sc_hd__o21a_1
XFILLER_65_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2040_ _2526_/A _2061_/B VGND VGND VPWR VPWR _2040_/X sky130_fd_sc_hd__or2_1
XFILLER_47_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2942_ _2961_/A VGND VGND VPWR VPWR _2956_/A sky130_fd_sc_hd__buf_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2873_ _3099_/B _2932_/B VGND VGND VPWR VPWR _2873_/X sky130_fd_sc_hd__or2_1
X_1824_ _2092_/C VGND VGND VPWR VPWR _2009_/B sky130_fd_sc_hd__clkbuf_2
X_1755_ _2832_/A VGND VGND VPWR VPWR _1755_/X sky130_fd_sc_hd__clkbuf_2
X_1686_ _2410_/A _2911_/A VGND VGND VPWR VPWR _1686_/Y sky130_fd_sc_hd__nor2_1
X_3356_ _2466_/Y _2463_/Y _3357_/S VGND VGND VPWR VPWR _3356_/X sky130_fd_sc_hd__mux2_1
X_3287_ _1784_/Y _1775_/Y _3351_/S VGND VGND VPWR VPWR _3287_/X sky130_fd_sc_hd__mux2_2
XFILLER_57_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2307_ _3058_/A _3094_/B VGND VGND VPWR VPWR _2307_/Y sky130_fd_sc_hd__nor2_1
X_2238_ _2202_/X _2605_/B _2237_/X VGND VGND VPWR VPWR _2238_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater275 _3347_/S VGND VGND VPWR VPWR _3380_/S sky130_fd_sc_hd__buf_6
X_2169_ _2426_/A VGND VGND VPWR VPWR _2390_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3210_ _2885_/Y _2881_/Y _3340_/S VGND VGND VPWR VPWR _3210_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3141_ _2638_/Y _2636_/Y _3340_/S VGND VGND VPWR VPWR _3141_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3072_ _3105_/A _3072_/B VGND VGND VPWR VPWR _3072_/X sky130_fd_sc_hd__or2_1
X_2023_ _2234_/A VGND VGND VPWR VPWR _2023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2925_ _2925_/A _2939_/A VGND VGND VPWR VPWR _2925_/X sky130_fd_sc_hd__or2_1
X_2856_ _2864_/A _2856_/B VGND VGND VPWR VPWR _2856_/Y sky130_fd_sc_hd__nor2_1
X_1807_ _2076_/A VGND VGND VPWR VPWR _2067_/A sky130_fd_sc_hd__clkbuf_2
X_2787_ _2794_/A _2787_/B VGND VGND VPWR VPWR _2787_/Y sky130_fd_sc_hd__nor2_1
X_1738_ _2239_/A _1732_/B _1709_/X VGND VGND VPWR VPWR _1740_/C sky130_fd_sc_hd__o21ai_2
X_1669_ _2042_/A _2268_/B _1605_/B _1951_/A VGND VGND VPWR VPWR _1673_/A sky130_fd_sc_hd__a31o_1
X_3408_ _3408_/CLK _3408_/D input1/X VGND VGND VPWR VPWR _3408_/Q sky130_fd_sc_hd__dfrtp_1
X_3339_ _2375_/Y _2369_/Y _3357_/S VGND VGND VPWR VPWR _3339_/X sky130_fd_sc_hd__mux2_2
XFILLER_26_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2710_ _1838_/B _2704_/X _2938_/B _2673_/X _2709_/X VGND VGND VPWR VPWR _2710_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2641_ _3099_/B _2641_/B VGND VGND VPWR VPWR _2641_/X sky130_fd_sc_hd__or2_1
X_2572_ _2572_/A VGND VGND VPWR VPWR _2577_/A sky130_fd_sc_hd__buf_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3124_ _3124_/A _3124_/B VGND VGND VPWR VPWR _3124_/X sky130_fd_sc_hd__or2_1
XFILLER_67_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3055_ _3052_/X _2828_/B _3053_/X _2593_/B _3054_/X VGND VGND VPWR VPWR _3055_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2006_ _2005_/X _1890_/A _1961_/X VGND VGND VPWR VPWR _2992_/B sky130_fd_sc_hd__a21oi_4
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2908_ _2674_/A _2901_/X _2872_/X _2672_/B _2907_/X VGND VGND VPWR VPWR _2908_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2839_ _2839_/A _2839_/B VGND VGND VPWR VPWR _2839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2624_ _3077_/B _2602_/X _2594_/X _2853_/B _2623_/X VGND VGND VPWR VPWR _2624_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput113 _3349_/X VGND VGND VPWR VPWR output_thermometer_o[221] sky130_fd_sc_hd__clkbuf_2
Xoutput124 _3298_/X VGND VGND VPWR VPWR output_thermometer_o[170] sky130_fd_sc_hd__clkbuf_2
Xoutput102 _3329_/X VGND VGND VPWR VPWR output_thermometer_o[201] sky130_fd_sc_hd__clkbuf_2
X_2555_ _2315_/X _3024_/B _2554_/X VGND VGND VPWR VPWR _2555_/Y sky130_fd_sc_hd__o21ai_1
Xoutput157 _3274_/X VGND VGND VPWR VPWR output_thermometer_o[146] sky130_fd_sc_hd__clkbuf_2
Xoutput135 _3140_/X VGND VGND VPWR VPWR output_thermometer_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput168 _3246_/X VGND VGND VPWR VPWR output_thermometer_o[118] sky130_fd_sc_hd__clkbuf_2
Xoutput146 _3217_/X VGND VGND VPWR VPWR output_thermometer_o[89] sky130_fd_sc_hd__clkbuf_2
Xoutput179 _3233_/X VGND VGND VPWR VPWR output_thermometer_o[105] sky130_fd_sc_hd__clkbuf_2
X_2486_ _2486_/A _2495_/B VGND VGND VPWR VPWR _2968_/B sky130_fd_sc_hd__or2_1
X_3107_ _3107_/A _3107_/B VGND VGND VPWR VPWR _3107_/Y sky130_fd_sc_hd__nor2_1
X_3038_ _3041_/A _3038_/B VGND VGND VPWR VPWR _3038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2340_ _2340_/A VGND VGND VPWR VPWR _3104_/B sky130_fd_sc_hd__inv_2
X_2271_ _2271_/A VGND VGND VPWR VPWR _2271_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1986_ _1951_/X _1982_/A _1961_/X VGND VGND VPWR VPWR _2985_/B sky130_fd_sc_hd__a21oi_4
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ _2607_/A VGND VGND VPWR VPWR _2607_/X sky130_fd_sc_hd__buf_2
X_2538_ _2538_/A VGND VGND VPWR VPWR _2538_/Y sky130_fd_sc_hd__inv_2
X_2469_ _2454_/X _2952_/B _1878_/B _2464_/X VGND VGND VPWR VPWR _2469_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ _1900_/A VGND VGND VPWR VPWR _1840_/X sky130_fd_sc_hd__buf_4
X_1771_ _1735_/X _2694_/B _1770_/X VGND VGND VPWR VPWR _1771_/Y sky130_fd_sc_hd__o21ai_1
X_3372_ _2536_/Y _2534_/Y _3374_/S VGND VGND VPWR VPWR _3372_/X sky130_fd_sc_hd__mux2_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2323_ _3099_/C VGND VGND VPWR VPWR _3054_/A sky130_fd_sc_hd__clkbuf_2
X_2254_ _2615_/B VGND VGND VPWR VPWR _2254_/Y sky130_fd_sc_hd__inv_2
X_2185_ _2185_/A VGND VGND VPWR VPWR _2185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1969_ _1981_/A _2310_/A VGND VGND VPWR VPWR _1970_/A sky130_fd_sc_hd__or2_2
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2941_ _2960_/A VGND VGND VPWR VPWR _2941_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2872_ _2960_/A VGND VGND VPWR VPWR _2872_/X sky130_fd_sc_hd__buf_2
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1823_ _3044_/A _1823_/B VGND VGND VPWR VPWR _2703_/B sky130_fd_sc_hd__nor2_4
X_1754_ _2185_/A _1756_/C VGND VGND VPWR VPWR _2431_/A sky130_fd_sc_hd__or2_2
X_1685_ _1689_/B VGND VGND VPWR VPWR _2911_/A sky130_fd_sc_hd__inv_2
X_3355_ _2461_/Y _2458_/Y _3383_/S VGND VGND VPWR VPWR _3355_/X sky130_fd_sc_hd__mux2_1
X_3286_ _1771_/Y _1765_/Y _3347_/S VGND VGND VPWR VPWR _3286_/X sky130_fd_sc_hd__mux2_4
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2306_ _2310_/A _2338_/A VGND VGND VPWR VPWR _3094_/B sky130_fd_sc_hd__nor2_2
X_2237_ _2315_/A _2839_/B _2206_/X _3064_/B VGND VGND VPWR VPWR _2237_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater276 _3382_/S VGND VGND VPWR VPWR _3347_/S sky130_fd_sc_hd__buf_6
X_2168_ _2168_/A _2168_/B VGND VGND VPWR VPWR _2426_/A sky130_fd_sc_hd__or2_1
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2099_ _1639_/X _2548_/A _2291_/A _1988_/A _2841_/A VGND VGND VPWR VPWR _2100_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3140_ _2635_/Y _2633_/Y _3342_/S VGND VGND VPWR VPWR _3140_/X sky130_fd_sc_hd__mux2_2
X_3071_ _3083_/A _3071_/B VGND VGND VPWR VPWR _3071_/Y sky130_fd_sc_hd__nor2_1
X_2022_ _2022_/A VGND VGND VPWR VPWR _2522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2924_ _2924_/A _2924_/B VGND VGND VPWR VPWR _2924_/Y sky130_fd_sc_hd__nor2_1
X_2855_ _2825_/X _3077_/B _2833_/X _2621_/B _2854_/X VGND VGND VPWR VPWR _2855_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1806_ _2157_/A VGND VGND VPWR VPWR _1806_/X sky130_fd_sc_hd__clkbuf_4
X_2786_ _2075_/B _2761_/X _3014_/B _2773_/X _2785_/X VGND VGND VPWR VPWR _2786_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1737_ _2030_/A VGND VGND VPWR VPWR _2239_/A sky130_fd_sc_hd__buf_2
X_1668_ _2092_/C _2157_/C VGND VGND VPWR VPWR _1951_/A sky130_fd_sc_hd__nor2_2
X_3407_ _3408_/CLK _3407_/D input1/X VGND VGND VPWR VPWR _3408_/D sky130_fd_sc_hd__dfrtp_1
X_1599_ _2113_/A VGND VGND VPWR VPWR _2092_/C sky130_fd_sc_hd__clkbuf_2
X_3338_ _2366_/Y _2360_/Y _3354_/S VGND VGND VPWR VPWR _3338_/X sky130_fd_sc_hd__mux2_2
XFILLER_65_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3269_ _3095_/Y _3093_/Y _3340_/S VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2640_ _2659_/A _2640_/B VGND VGND VPWR VPWR _2640_/Y sky130_fd_sc_hd__nor2_1
X_2571_ input2/X _3408_/D _2165_/B _2401_/A VGND VGND VPWR VPWR _2571_/X sky130_fd_sc_hd__a31o_1
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3123_ _3126_/A _3123_/B VGND VGND VPWR VPWR _3123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3054_ _3054_/A _3054_/B VGND VGND VPWR VPWR _3054_/X sky130_fd_sc_hd__or2_1
X_2005_ _2067_/A VGND VGND VPWR VPWR _2005_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2907_ _2907_/A _2922_/B VGND VGND VPWR VPWR _2907_/X sky130_fd_sc_hd__or2_1
X_2838_ _2087_/X _2600_/B _1797_/X _3062_/B _2837_/X VGND VGND VPWR VPWR _2838_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2769_ _2776_/A _2769_/B VGND VGND VPWR VPWR _2769_/Y sky130_fd_sc_hd__nor2_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2623_ _3081_/B _2641_/B VGND VGND VPWR VPWR _2623_/X sky130_fd_sc_hd__or2_1
Xoutput114 _3224_/X VGND VGND VPWR VPWR output_thermometer_o[96] sky130_fd_sc_hd__clkbuf_2
Xoutput125 _3288_/X VGND VGND VPWR VPWR output_thermometer_o[160] sky130_fd_sc_hd__clkbuf_2
Xoutput103 _3311_/X VGND VGND VPWR VPWR output_thermometer_o[183] sky130_fd_sc_hd__clkbuf_2
X_2554_ _2794_/B _2294_/X _3025_/B _2549_/X VGND VGND VPWR VPWR _2554_/X sky130_fd_sc_hd__o22a_1
Xoutput158 _3353_/X VGND VGND VPWR VPWR output_thermometer_o[225] sky130_fd_sc_hd__clkbuf_2
Xoutput147 _3303_/X VGND VGND VPWR VPWR output_thermometer_o[175] sky130_fd_sc_hd__clkbuf_2
Xoutput136 _3261_/X VGND VGND VPWR VPWR output_thermometer_o[133] sky130_fd_sc_hd__clkbuf_2
Xoutput169 _3319_/X VGND VGND VPWR VPWR output_thermometer_o[191] sky130_fd_sc_hd__clkbuf_2
X_2485_ _2730_/B _2483_/X _2484_/X VGND VGND VPWR VPWR _2485_/Y sky130_fd_sc_hd__o21ai_1
X_3106_ _1777_/X _2645_/B _2097_/X _2343_/Y _3105_/X VGND VGND VPWR VPWR _3106_/Y
+ sky130_fd_sc_hd__o221ai_2
X_3037_ _2806_/A _2607_/X _3032_/X _2805_/B _3036_/X VGND VGND VPWR VPWR _3037_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2270_ _1769_/B _2266_/A _1631_/B _1900_/A VGND VGND VPWR VPWR _2271_/A sky130_fd_sc_hd__a31o_1
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1985_ _1996_/A _1985_/B VGND VGND VPWR VPWR _1985_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2606_ _2606_/A VGND VGND VPWR VPWR _2606_/X sky130_fd_sc_hd__clkbuf_2
X_2537_ _2537_/A _2785_/B VGND VGND VPWR VPWR _2538_/A sky130_fd_sc_hd__or2_2
X_2468_ _2953_/B VGND VGND VPWR VPWR _2468_/Y sky130_fd_sc_hd__inv_2
X_2399_ _3124_/B VGND VGND VPWR VPWR _2399_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1770_ _1708_/X _2434_/A _1755_/X _2928_/B VGND VGND VPWR VPWR _1770_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3371_ _2533_/Y _2530_/Y _3374_/S VGND VGND VPWR VPWR _3371_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2322_ _2322_/A VGND VGND VPWR VPWR _3102_/B sky130_fd_sc_hd__inv_2
X_2253_ _2398_/A _3072_/B VGND VGND VPWR VPWR _2615_/B sky130_fd_sc_hd__or2_1
X_2184_ _2184_/A VGND VGND VPWR VPWR _2184_/X sky130_fd_sc_hd__buf_2
X_1968_ _1968_/A VGND VGND VPWR VPWR _2310_/A sky130_fd_sc_hd__clkinv_4
X_1899_ _1938_/A _1899_/B VGND VGND VPWR VPWR _1899_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2940_ _3001_/A VGND VGND VPWR VPWR _2940_/X sky130_fd_sc_hd__clkbuf_2
X_2871_ _2886_/A _2871_/B VGND VGND VPWR VPWR _2871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1822_ _2242_/A VGND VGND VPWR VPWR _3044_/A sky130_fd_sc_hd__buf_2
X_1753_ _2239_/A _1747_/B _1709_/X VGND VGND VPWR VPWR _1756_/C sky130_fd_sc_hd__o21ai_1
X_1684_ _1684_/A _1684_/B _1747_/C VGND VGND VPWR VPWR _1689_/B sky130_fd_sc_hd__or3_4
X_3354_ _2456_/Y _2453_/Y _3354_/S VGND VGND VPWR VPWR _3354_/X sky130_fd_sc_hd__mux2_2
X_3285_ _1758_/Y _1749_/Y _3347_/S VGND VGND VPWR VPWR _3285_/X sky130_fd_sc_hd__mux2_4
X_2305_ _2202_/X _2633_/B _2304_/X VGND VGND VPWR VPWR _2305_/Y sky130_fd_sc_hd__o21ai_1
X_2236_ _2236_/A VGND VGND VPWR VPWR _3064_/B sky130_fd_sc_hd__inv_2
XFILLER_57_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater277 _3342_/S VGND VGND VPWR VPWR _3382_/S sky130_fd_sc_hd__buf_8
X_2167_ _2301_/C _1789_/X _2851_/A _2166_/X VGND VGND VPWR VPWR _2167_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2098_ _2889_/A VGND VGND VPWR VPWR _3027_/A sky130_fd_sc_hd__buf_2
XFILLER_21_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3070_ _3052_/X _2845_/B _3053_/X _2610_/B _3069_/X VGND VGND VPWR VPWR _3070_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2021_ _2195_/A VGND VGND VPWR VPWR _2022_/A sky130_fd_sc_hd__inv_2
XFILLER_47_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2923_ _1740_/C _2920_/X _2921_/X _2688_/B _2922_/X VGND VGND VPWR VPWR _2923_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2854_ _3081_/B _2854_/B VGND VGND VPWR VPWR _2854_/X sky130_fd_sc_hd__or2_1
X_2785_ _2785_/A _2785_/B _2785_/C VGND VGND VPWR VPWR _2785_/X sky130_fd_sc_hd__or3_1
X_1805_ _2113_/A VGND VGND VPWR VPWR _2157_/A sky130_fd_sc_hd__buf_2
X_1736_ _2089_/A _1736_/B VGND VGND VPWR VPWR _2688_/B sky130_fd_sc_hd__nor2_4
X_1667_ _2018_/A VGND VGND VPWR VPWR _2157_/C sky130_fd_sc_hd__clkbuf_2
X_1598_ _1588_/Y _1642_/A _2178_/A _2932_/A VGND VGND VPWR VPWR _2113_/A sky130_fd_sc_hd__a31o_2
X_3406_ _3408_/CLK _3406_/D input1/X VGND VGND VPWR VPWR _3407_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_58_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3337_ _2357_/Y _2350_/Y _3357_/S VGND VGND VPWR VPWR _3337_/X sky130_fd_sc_hd__mux2_1
X_3268_ _3092_/Y _3090_/Y _3354_/S VGND VGND VPWR VPWR _3268_/X sky130_fd_sc_hd__mux2_2
X_2219_ _2219_/A _2219_/B VGND VGND VPWR VPWR _3062_/B sky130_fd_sc_hd__nand2_2
X_3199_ _2850_/X _2848_/Y _3351_/S VGND VGND VPWR VPWR _3199_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2570_ _1653_/X _3041_/B _2569_/X VGND VGND VPWR VPWR _2570_/Y sky130_fd_sc_hd__o21ai_1
X_3122_ _1653_/X _2663_/B _3121_/X VGND VGND VPWR VPWR _3122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3053_ _3098_/A VGND VGND VPWR VPWR _3053_/X sky130_fd_sc_hd__clkbuf_2
X_2004_ _2056_/A _2004_/B VGND VGND VPWR VPWR _2004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2906_ _3004_/A VGND VGND VPWR VPWR _2922_/B sky130_fd_sc_hd__clkbuf_2
X_2837_ _2837_/A _3060_/B _2879_/C VGND VGND VPWR VPWR _2837_/X sky130_fd_sc_hd__or3_2
X_2768_ _2522_/A _2763_/X _2996_/B _2753_/X _2767_/X VGND VGND VPWR VPWR _2768_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1719_ _1721_/B VGND VGND VPWR VPWR _2917_/A sky130_fd_sc_hd__inv_2
X_2699_ _2440_/A _2653_/X _2931_/B _2673_/X _2698_/X VGND VGND VPWR VPWR _2699_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2622_ _2792_/B VGND VGND VPWR VPWR _2641_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput104 _3365_/X VGND VGND VPWR VPWR output_thermometer_o[237] sky130_fd_sc_hd__clkbuf_2
X_2553_ _2565_/A _2795_/A VGND VGND VPWR VPWR _2553_/Y sky130_fd_sc_hd__nor2_1
Xoutput115 _3202_/X VGND VGND VPWR VPWR output_thermometer_o[74] sky130_fd_sc_hd__clkbuf_2
Xoutput126 _3228_/X VGND VGND VPWR VPWR output_thermometer_o[100] sky130_fd_sc_hd__clkbuf_2
Xoutput137 _3295_/X VGND VGND VPWR VPWR output_thermometer_o[167] sky130_fd_sc_hd__clkbuf_2
Xoutput159 _3236_/X VGND VGND VPWR VPWR output_thermometer_o[108] sky130_fd_sc_hd__clkbuf_2
Xoutput148 _3212_/X VGND VGND VPWR VPWR output_thermometer_o[84] sky130_fd_sc_hd__clkbuf_2
X_2484_ _2478_/X _2964_/B _1912_/B _2464_/X VGND VGND VPWR VPWR _2484_/X sky130_fd_sc_hd__o22a_1
X_3105_ _3105_/A _3105_/B VGND VGND VPWR VPWR _3105_/X sky130_fd_sc_hd__or2_1
X_3036_ _3042_/A _3036_/B VGND VGND VPWR VPWR _3036_/X sky130_fd_sc_hd__or2_1
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1984_ _1987_/B VGND VGND VPWR VPWR _1985_/B sky130_fd_sc_hd__inv_2
XFILLER_60_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2605_ _2610_/A _2605_/B VGND VGND VPWR VPWR _2605_/Y sky130_fd_sc_hd__nor2_1
X_2536_ _2776_/B _2527_/X _2535_/X VGND VGND VPWR VPWR _2536_/Y sky130_fd_sc_hd__o21ai_1
X_2467_ _2467_/A _2471_/B VGND VGND VPWR VPWR _2953_/B sky130_fd_sc_hd__or2_2
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2398_ _2398_/A _2398_/B VGND VGND VPWR VPWR _3124_/B sky130_fd_sc_hd__or2_2
X_3019_ _3019_/A _3019_/B VGND VGND VPWR VPWR _3019_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3370_ _2529_/Y _2526_/Y _3370_/S VGND VGND VPWR VPWR _3370_/X sky130_fd_sc_hd__mux2_2
X_2321_ _2265_/A _2265_/B _2161_/Y VGND VGND VPWR VPWR _2322_/A sky130_fd_sc_hd__o21ai_2
XFILLER_2_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2252_ _2265_/A _2252_/B VGND VGND VPWR VPWR _3072_/B sky130_fd_sc_hd__nor2_2
X_2183_ _2233_/A VGND VGND VPWR VPWR _2184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ _1913_/X _2977_/B _1963_/X _2746_/B _1966_/X VGND VGND VPWR VPWR _1967_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1898_ _1903_/B VGND VGND VPWR VPWR _1899_/B sky130_fd_sc_hd__inv_2
XFILLER_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2519_ _2501_/X _2992_/B _2004_/B _2511_/X VGND VGND VPWR VPWR _2519_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2870_ _2857_/X _3093_/B _2833_/X _2636_/B _2869_/X VGND VGND VPWR VPWR _2870_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1821_ _1820_/X _1811_/A _1779_/A VGND VGND VPWR VPWR _2935_/B sky130_fd_sc_hd__a21oi_4
X_1752_ _2232_/A _1752_/B VGND VGND VPWR VPWR _2691_/B sky130_fd_sc_hd__nor2_2
X_1683_ _1683_/A VGND VGND VPWR VPWR _1747_/C sky130_fd_sc_hd__clkbuf_2
X_3353_ _2449_/Y _2447_/Y _3354_/S VGND VGND VPWR VPWR _3353_/X sky130_fd_sc_hd__mux2_1
X_3284_ _1742_/Y _1734_/Y _3347_/S VGND VGND VPWR VPWR _3284_/X sky130_fd_sc_hd__mux2_2
X_2304_ _2246_/X _2864_/B _2097_/X _3090_/A VGND VGND VPWR VPWR _2304_/X sky130_fd_sc_hd__o22a_1
X_2235_ _2233_/X _2229_/B _2234_/X VGND VGND VPWR VPWR _2839_/B sky130_fd_sc_hd__o21a_1
X_2166_ _2166_/A VGND VGND VPWR VPWR _2166_/X sky130_fd_sc_hd__buf_1
Xrepeater278 _3330_/S VGND VGND VPWR VPWR _3340_/S sky130_fd_sc_hd__buf_8
X_2097_ _2727_/A VGND VGND VPWR VPWR _2097_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2999_ _2522_/A _2994_/X _2997_/X _2765_/B _2998_/X VGND VGND VPWR VPWR _2999_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2020_ _2103_/A VGND VGND VPWR VPWR _2020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2922_ _2922_/A _2922_/B VGND VGND VPWR VPWR _2922_/X sky130_fd_sc_hd__or2_1
XFILLER_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2853_ _2864_/A _2853_/B VGND VGND VPWR VPWR _2853_/Y sky130_fd_sc_hd__nor2_1
X_2784_ _2794_/A _2784_/B VGND VGND VPWR VPWR _2784_/Y sky130_fd_sc_hd__nor2_1
X_1804_ _2568_/A VGND VGND VPWR VPWR _1878_/A sky130_fd_sc_hd__clkbuf_2
X_1735_ _2131_/A VGND VGND VPWR VPWR _1735_/X sky130_fd_sc_hd__clkbuf_2
X_1666_ _1683_/A VGND VGND VPWR VPWR _2018_/A sky130_fd_sc_hd__inv_2
X_1597_ _1773_/B VGND VGND VPWR VPWR _2932_/A sky130_fd_sc_hd__inv_2
X_3405_ _3408_/CLK _3405_/D input1/X VGND VGND VPWR VPWR _3406_/D sky130_fd_sc_hd__dfrtp_1
X_3336_ _2346_/Y _2339_/Y _3351_/S VGND VGND VPWR VPWR _3336_/X sky130_fd_sc_hd__mux2_2
X_3267_ _3089_/Y _3087_/Y _3340_/S VGND VGND VPWR VPWR _3267_/X sky130_fd_sc_hd__mux2_1
X_2218_ _2397_/A _2221_/B VGND VGND VPWR VPWR _2219_/B sky130_fd_sc_hd__or2_2
X_3198_ _2847_/Y _2845_/Y _3330_/S VGND VGND VPWR VPWR _3198_/X sky130_fd_sc_hd__mux2_2
X_2149_ _2149_/A _2149_/B _2157_/C VGND VGND VPWR VPWR _2809_/A sky130_fd_sc_hd__or3_4
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3121_ _1818_/A _2894_/B _1610_/X _2388_/A VGND VGND VPWR VPWR _3121_/X sky130_fd_sc_hd__o22a_1
XFILLER_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3052_ _3097_/A VGND VGND VPWR VPWR _3052_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2003_ _2007_/B VGND VGND VPWR VPWR _2004_/B sky130_fd_sc_hd__inv_2
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2905_ _2905_/A _2905_/B VGND VGND VPWR VPWR _2905_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2836_ _2839_/A _2836_/B VGND VGND VPWR VPWR _2836_/Y sky130_fd_sc_hd__nor2_1
X_2767_ _2998_/B _2782_/B VGND VGND VPWR VPWR _2767_/X sky130_fd_sc_hd__or2_1
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1718_ _1763_/A _1718_/B _1747_/C VGND VGND VPWR VPWR _1721_/B sky130_fd_sc_hd__or3_4
X_2698_ _2932_/A _2792_/B VGND VGND VPWR VPWR _2698_/X sky130_fd_sc_hd__or2_1
X_1649_ _1639_/X _2548_/A _2391_/A VGND VGND VPWR VPWR _1658_/B sky130_fd_sc_hd__o21ai_4
X_3319_ _2167_/X _2161_/Y _3351_/S VGND VGND VPWR VPWR _3319_/X sky130_fd_sc_hd__mux2_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2621_ _2636_/A _2621_/B VGND VGND VPWR VPWR _2621_/Y sky130_fd_sc_hd__nor2_1
X_2552_ _3110_/A VGND VGND VPWR VPWR _2565_/A sky130_fd_sc_hd__clkbuf_2
Xoutput105 _3172_/X VGND VGND VPWR VPWR output_thermometer_o[44] sky130_fd_sc_hd__clkbuf_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput116 _3335_/X VGND VGND VPWR VPWR output_thermometer_o[207] sky130_fd_sc_hd__clkbuf_2
Xoutput138 _3332_/X VGND VGND VPWR VPWR output_thermometer_o[204] sky130_fd_sc_hd__clkbuf_2
Xoutput127 _3213_/X VGND VGND VPWR VPWR output_thermometer_o[85] sky130_fd_sc_hd__clkbuf_2
Xoutput149 _3378_/X VGND VGND VPWR VPWR output_thermometer_o[250] sky130_fd_sc_hd__clkbuf_2
X_2483_ _2527_/A VGND VGND VPWR VPWR _2483_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3104_ _3107_/A _3104_/B VGND VGND VPWR VPWR _3104_/Y sky130_fd_sc_hd__nor2_1
X_3035_ _3041_/A _3035_/B VGND VGND VPWR VPWR _3035_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2819_ _3032_/A _2939_/A VGND VGND VPWR VPWR _2820_/A sky130_fd_sc_hd__nand2_2
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1983_ _1931_/X _2509_/A _1935_/X VGND VGND VPWR VPWR _1987_/B sky130_fd_sc_hd__o21ai_2
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2604_ _3060_/B _2602_/X _2594_/X _2836_/B _2603_/X VGND VGND VPWR VPWR _2604_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2535_ _2523_/X _3008_/B _3009_/B _2531_/X VGND VGND VPWR VPWR _2535_/X sky130_fd_sc_hd__o22a_1
X_2466_ _2714_/B _2459_/X _2465_/X VGND VGND VPWR VPWR _2466_/Y sky130_fd_sc_hd__o21ai_1
X_2397_ _2397_/A _2400_/B VGND VGND VPWR VPWR _2398_/B sky130_fd_sc_hd__nor2_2
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3018_ _3024_/A _3018_/B VGND VGND VPWR VPWR _3018_/Y sky130_fd_sc_hd__nor2_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2320_ _2315_/X _2871_/B _2319_/X VGND VGND VPWR VPWR _2320_/Y sky130_fd_sc_hd__o21ai_1
X_2251_ _2202_/X _2610_/B _2250_/X VGND VGND VPWR VPWR _2251_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2182_ _2290_/A _3049_/B VGND VGND VPWR VPWR _2182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1966_ _1978_/A _2499_/A _2071_/C VGND VGND VPWR VPWR _1966_/X sky130_fd_sc_hd__or3_2
X_1897_ _1871_/X _2476_/A _1875_/X VGND VGND VPWR VPWR _1903_/B sky130_fd_sc_hd__o21ai_2
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2518_ _2993_/B VGND VGND VPWR VPWR _2518_/Y sky130_fd_sc_hd__inv_2
X_2449_ _2703_/B _2428_/X _2448_/X VGND VGND VPWR VPWR _2449_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1820_ _1890_/A VGND VGND VPWR VPWR _1820_/X sky130_fd_sc_hd__buf_4
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _2242_/A VGND VGND VPWR VPWR _2232_/A sky130_fd_sc_hd__buf_4
X_1682_ _2114_/B VGND VGND VPWR VPWR _1684_/B sky130_fd_sc_hd__inv_2
X_3352_ _2445_/Y _2443_/Y _3382_/S VGND VGND VPWR VPWR _3352_/X sky130_fd_sc_hd__mux2_1
X_2303_ _2082_/A _2184_/A _2499_/A _2158_/A VGND VGND VPWR VPWR _3090_/A sky130_fd_sc_hd__a31o_2
X_3283_ _1727_/Y _1720_/Y _3347_/S VGND VGND VPWR VPWR _3283_/X sky130_fd_sc_hd__mux2_2
X_2234_ _2234_/A VGND VGND VPWR VPWR _2234_/X sky130_fd_sc_hd__clkbuf_2
X_2165_ _2242_/A _2165_/B VGND VGND VPWR VPWR _2166_/A sky130_fd_sc_hd__or2_1
Xrepeater279 _3342_/S VGND VGND VPWR VPWR _3330_/S sky130_fd_sc_hd__buf_8
X_2096_ _2401_/A _2096_/B VGND VGND VPWR VPWR _2790_/B sky130_fd_sc_hd__nor2_4
XFILLER_53_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2998_ _3001_/A _2998_/B VGND VGND VPWR VPWR _2998_/X sky130_fd_sc_hd__or2_1
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1949_ _1953_/B VGND VGND VPWR VPWR _1950_/B sky130_fd_sc_hd__inv_2
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2921_ _2960_/A VGND VGND VPWR VPWR _2921_/X sky130_fd_sc_hd__clkbuf_4
X_2852_ _2301_/C _1789_/X _3074_/B _2821_/B _2851_/Y VGND VGND VPWR VPWR _2852_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1803_ _1789_/X _1794_/Y _1797_/X _1799_/Y _1802_/X VGND VGND VPWR VPWR _1803_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2783_ _1789_/X _2538_/A _3011_/B _2773_/X _2782_/X VGND VGND VPWR VPWR _2783_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1734_ _1786_/A _2922_/A VGND VGND VPWR VPWR _1734_/Y sky130_fd_sc_hd__nor2_1
X_1665_ _1744_/A VGND VGND VPWR VPWR _2268_/B sky130_fd_sc_hd__clkbuf_2
X_3404_ _3404_/CLK _3404_/D input1/X VGND VGND VPWR VPWR _3405_/D sky130_fd_sc_hd__dfrtp_1
X_1596_ _1860_/A _1570_/A _2101_/A VGND VGND VPWR VPWR _1773_/B sky130_fd_sc_hd__o21ai_1
X_3335_ _2337_/Y _3102_/B _3354_/S VGND VGND VPWR VPWR _3335_/X sky130_fd_sc_hd__mux2_2
X_3266_ _3085_/Y _3083_/Y _3330_/S VGND VGND VPWR VPWR _3266_/X sky130_fd_sc_hd__mux2_1
X_2217_ _2212_/X _2831_/B _2216_/X VGND VGND VPWR VPWR _2217_/Y sky130_fd_sc_hd__o21ai_1
X_3197_ _2843_/Y _2839_/Y _3342_/S VGND VGND VPWR VPWR _3197_/X sky130_fd_sc_hd__mux2_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2148_ _2156_/A _2148_/B VGND VGND VPWR VPWR _2808_/B sky130_fd_sc_hd__nor2_2
XFILLER_53_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2079_ _2245_/A VGND VGND VPWR VPWR _3098_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3120_ _3120_/A VGND VGND VPWR VPWR _3120_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3051_ _3064_/A _3051_/B VGND VGND VPWR VPWR _3051_/Y sky130_fd_sc_hd__nor2_1
X_2002_ _1639_/X _1806_/X _2291_/A VGND VGND VPWR VPWR _2007_/B sky130_fd_sc_hd__o21ai_4
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2904_ _1632_/C _2901_/X _2669_/B _1818_/X _2903_/X VGND VGND VPWR VPWR _2904_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_31_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2835_ _2825_/X _3056_/B _2833_/X _2597_/B _2834_/X VGND VGND VPWR VPWR _2835_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2766_ _2766_/A VGND VGND VPWR VPWR _2782_/B sky130_fd_sc_hd__buf_1
X_1717_ _2133_/B VGND VGND VPWR VPWR _1718_/B sky130_fd_sc_hd__inv_2
X_2697_ _2931_/A _2697_/B VGND VGND VPWR VPWR _2697_/Y sky130_fd_sc_hd__nor2_1
X_1648_ _1648_/A VGND VGND VPWR VPWR _2391_/A sky130_fd_sc_hd__buf_2
X_3318_ _2160_/Y _2155_/Y _3382_/S VGND VGND VPWR VPWR _3318_/X sky130_fd_sc_hd__mux2_2
X_1579_ _2245_/A VGND VGND VPWR VPWR _2523_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3249_ _3026_/Y _3024_/Y _3381_/S VGND VGND VPWR VPWR _3249_/X sky130_fd_sc_hd__mux2_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ _2662_/A VGND VGND VPWR VPWR _2636_/A sky130_fd_sc_hd__clkbuf_2
X_2551_ _2790_/B _2545_/X _2550_/X VGND VGND VPWR VPWR _2551_/Y sky130_fd_sc_hd__o21ai_1
Xoutput106 _3262_/X VGND VGND VPWR VPWR output_thermometer_o[134] sky130_fd_sc_hd__clkbuf_2
Xoutput117 _3255_/X VGND VGND VPWR VPWR output_thermometer_o[127] sky130_fd_sc_hd__clkbuf_2
Xoutput139 _3350_/X VGND VGND VPWR VPWR output_thermometer_o[222] sky130_fd_sc_hd__clkbuf_2
Xoutput128 _3320_/X VGND VGND VPWR VPWR output_thermometer_o[192] sky130_fd_sc_hd__clkbuf_2
X_2482_ _2965_/B VGND VGND VPWR VPWR _2482_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3103_ _2577_/A _2335_/A _3102_/X _2851_/A _2617_/B VGND VGND VPWR VPWR _3103_/X
+ sky130_fd_sc_hd__a32o_1
X_3034_ _2803_/A _2607_/X _3032_/X _2802_/B _3033_/X VGND VGND VPWR VPWR _3034_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2818_ _3004_/A VGND VGND VPWR VPWR _2939_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2749_ _2756_/A _2749_/B VGND VGND VPWR VPWR _2749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1982_ _1982_/A VGND VGND VPWR VPWR _2509_/A sky130_fd_sc_hd__inv_2
X_2603_ _2705_/A _3062_/B VGND VGND VPWR VPWR _2603_/X sky130_fd_sc_hd__or2_1
X_2534_ _2534_/A _2548_/B VGND VGND VPWR VPWR _2534_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2465_ _2454_/X _2948_/B _1865_/B _2464_/X VGND VGND VPWR VPWR _2465_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2396_ _2315_/X _2894_/B _2395_/X VGND VGND VPWR VPWR _2396_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3017_ _2857_/A _2075_/B _3015_/X _2784_/B _3016_/Y VGND VGND VPWR VPWR _3017_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2250_ _2246_/X _2845_/B _2248_/X _3068_/B VGND VGND VPWR VPWR _2250_/X sky130_fd_sc_hd__o22a_1
X_2181_ _2195_/A _2289_/B VGND VGND VPWR VPWR _3049_/B sky130_fd_sc_hd__nor2_2
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1965_ _2082_/C VGND VGND VPWR VPWR _2071_/C sky130_fd_sc_hd__buf_1
X_1896_ _2252_/B VGND VGND VPWR VPWR _2476_/A sky130_fd_sc_hd__inv_2
X_2517_ _2756_/B _2506_/X _2516_/X VGND VGND VPWR VPWR _2517_/Y sky130_fd_sc_hd__o21ai_1
X_2448_ _2422_/X _2935_/B _1816_/B _2436_/X VGND VGND VPWR VPWR _2448_/X sky130_fd_sc_hd__o22a_1
X_2379_ _2347_/X _2058_/A _1648_/A VGND VGND VPWR VPWR _2383_/A sky130_fd_sc_hd__o21ai_4
XFILLER_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1750_ _2333_/A VGND VGND VPWR VPWR _2242_/A sky130_fd_sc_hd__buf_2
X_1681_ _2076_/A _1920_/A VGND VGND VPWR VPWR _2114_/B sky130_fd_sc_hd__nand2_4
X_3351_ _2441_/Y _2101_/Y _3351_/S VGND VGND VPWR VPWR _3351_/X sky130_fd_sc_hd__mux2_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2302_ _2233_/X _2299_/B _2142_/A VGND VGND VPWR VPWR _2864_/B sky130_fd_sc_hd__o21a_1
X_3282_ _1714_/Y _1706_/Y _3346_/S VGND VGND VPWR VPWR _3282_/X sky130_fd_sc_hd__mux2_2
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2233_ _2233_/A VGND VGND VPWR VPWR _2233_/X sky130_fd_sc_hd__clkbuf_2
X_2164_ _3019_/A VGND VGND VPWR VPWR _2851_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2095_ _2109_/A _2095_/B VGND VGND VPWR VPWR _2095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2997_ _3032_/A VGND VGND VPWR VPWR _2997_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1948_ _1931_/X _2495_/A _1935_/X VGND VGND VPWR VPWR _1953_/B sky130_fd_sc_hd__o21ai_2
X_1879_ _1820_/X _2231_/B _1840_/X VGND VGND VPWR VPWR _2952_/B sky130_fd_sc_hd__a21oi_4
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2920_ _2920_/A VGND VGND VPWR VPWR _2920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2851_ _2851_/A _2851_/B VGND VGND VPWR VPWR _2851_/Y sky130_fd_sc_hd__nand2_1
X_1802_ _1802_/A VGND VGND VPWR VPWR _1802_/X sky130_fd_sc_hd__clkbuf_2
X_2782_ _3012_/B _2782_/B VGND VGND VPWR VPWR _2782_/X sky130_fd_sc_hd__or2_1
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1733_ _1736_/B VGND VGND VPWR VPWR _2922_/A sky130_fd_sc_hd__inv_2
X_1664_ _1664_/A VGND VGND VPWR VPWR _1744_/A sky130_fd_sc_hd__clkbuf_2
X_3403_ _3404_/CLK _3403_/D input1/X VGND VGND VPWR VPWR _3404_/D sky130_fd_sc_hd__dfrtp_1
X_1595_ _2178_/A VGND VGND VPWR VPWR _2101_/A sky130_fd_sc_hd__inv_2
X_3334_ _2320_/Y _2314_/Y _3340_/S VGND VGND VPWR VPWR _3334_/X sky130_fd_sc_hd__mux2_2
X_3265_ _3082_/Y _3077_/Y _3330_/S VGND VGND VPWR VPWR _3265_/X sky130_fd_sc_hd__mux2_1
X_2216_ _2188_/X _3056_/B _2606_/A _2597_/B VGND VGND VPWR VPWR _2216_/X sky130_fd_sc_hd__o22a_1
X_3196_ _2838_/Y _2836_/Y _3346_/S VGND VGND VPWR VPWR _3196_/X sky130_fd_sc_hd__mux2_2
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2147_ _2155_/A _3039_/B VGND VGND VPWR VPWR _2147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2078_ _1890_/A _2400_/B _1900_/A VGND VGND VPWR VPWR _3014_/B sky130_fd_sc_hd__a21oi_4
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3050_ _2882_/X _2823_/B _2080_/X _2588_/B _3049_/X VGND VGND VPWR VPWR _3050_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2001_ _3047_/A VGND VGND VPWR VPWR _2056_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2903_ _3126_/B _3042_/A VGND VGND VPWR VPWR _2903_/X sky130_fd_sc_hd__or2_1
XFILLER_31_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2834_ _3058_/B _2854_/B VGND VGND VPWR VPWR _2834_/X sky130_fd_sc_hd__or2_1
X_2765_ _2776_/A _2765_/B VGND VGND VPWR VPWR _2765_/Y sky130_fd_sc_hd__nor2_1
X_2696_ _2928_/B _2682_/X _2695_/X VGND VGND VPWR VPWR _2696_/Y sky130_fd_sc_hd__o21ai_1
X_1716_ _1761_/A _1945_/A VGND VGND VPWR VPWR _2133_/B sky130_fd_sc_hd__or2_4
X_1647_ _2400_/A VGND VGND VPWR VPWR _1648_/A sky130_fd_sc_hd__inv_2
X_3317_ _2152_/Y _2147_/Y _3380_/S VGND VGND VPWR VPWR _3317_/X sky130_fd_sc_hd__mux2_1
X_1578_ _2168_/B _2993_/A VGND VGND VPWR VPWR _2245_/A sky130_fd_sc_hd__or2_2
X_3248_ _3023_/Y _3021_/Y _3382_/S VGND VGND VPWR VPWR _3248_/X sky130_fd_sc_hd__mux2_2
X_3179_ _2775_/Y _2772_/Y _3370_/S VGND VGND VPWR VPWR _3179_/X sky130_fd_sc_hd__mux2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ _1653_/A _2100_/B _2095_/B _2549_/X VGND VGND VPWR VPWR _2550_/X sky130_fd_sc_hd__o22a_1
Xoutput107 _3163_/X VGND VGND VPWR VPWR output_thermometer_o[35] sky130_fd_sc_hd__clkbuf_2
Xoutput129 _3176_/X VGND VGND VPWR VPWR output_thermometer_o[48] sky130_fd_sc_hd__clkbuf_2
X_2481_ _2481_/A _2495_/B VGND VGND VPWR VPWR _2965_/B sky130_fd_sc_hd__or2_1
Xoutput118 _3148_/X VGND VGND VPWR VPWR output_thermometer_o[20] sky130_fd_sc_hd__clkbuf_2
X_3102_ _3102_/A _3102_/B VGND VGND VPWR VPWR _3102_/X sky130_fd_sc_hd__or2_1
X_3033_ _3042_/A _3033_/B VGND VGND VPWR VPWR _3033_/X sky130_fd_sc_hd__or2_1
XFILLER_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2817_ _2817_/A VGND VGND VPWR VPWR _3032_/A sky130_fd_sc_hd__clkbuf_2
X_2748_ _1960_/B _2743_/X _2977_/B _2734_/X _2747_/X VGND VGND VPWR VPWR _2748_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2679_ _2889_/A VGND VGND VPWR VPWR _2759_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1981_ _1981_/A _2318_/A VGND VGND VPWR VPWR _1982_/A sky130_fd_sc_hd__or2_2
X_2602_ _2723_/A VGND VGND VPWR VPWR _2602_/X sky130_fd_sc_hd__buf_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2533_ _2772_/B _2527_/X _2532_/X VGND VGND VPWR VPWR _2533_/Y sky130_fd_sc_hd__o21ai_1
X_2464_ _2531_/A VGND VGND VPWR VPWR _2464_/X sky130_fd_sc_hd__clkbuf_2
X_2395_ _2390_/X _2663_/B _2393_/X _3120_/A VGND VGND VPWR VPWR _2395_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3016_ _3019_/A _3016_/B VGND VGND VPWR VPWR _3016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ _2338_/A VGND VGND VPWR VPWR _2289_/B sky130_fd_sc_hd__buf_2
XFILLER_65_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1964_ _1964_/A _1964_/B VGND VGND VPWR VPWR _2746_/B sky130_fd_sc_hd__nor2_2
X_1895_ _1907_/A _2257_/A VGND VGND VPWR VPWR _2252_/B sky130_fd_sc_hd__or2_4
X_2516_ _2501_/X _2989_/B _1996_/B _2511_/X VGND VGND VPWR VPWR _2516_/X sky130_fd_sc_hd__o22a_1
X_2447_ _2936_/B VGND VGND VPWR VPWR _2447_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2378_ _3118_/B VGND VGND VPWR VPWR _2378_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1680_ _3385_/Q _1809_/B _1808_/B _1744_/A VGND VGND VPWR VPWR _1920_/A sky130_fd_sc_hd__o31a_1
X_3350_ _2438_/Y _2434_/Y _3380_/S VGND VGND VPWR VPWR _3350_/X sky130_fd_sc_hd__mux2_1
X_2301_ _2301_/A _2499_/A _2301_/C VGND VGND VPWR VPWR _2633_/B sky130_fd_sc_hd__and3_2
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3281_ _1697_/Y _1686_/Y _3347_/S VGND VGND VPWR VPWR _3281_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2232_ _2232_/A _2236_/A VGND VGND VPWR VPWR _2605_/B sky130_fd_sc_hd__nor2_2
X_2163_ _2961_/A VGND VGND VPWR VPWR _3019_/A sky130_fd_sc_hd__inv_2
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2094_ _2096_/B VGND VGND VPWR VPWR _2095_/B sky130_fd_sc_hd__inv_2
XFILLER_53_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2996_ _3003_/A _2996_/B VGND VGND VPWR VPWR _2996_/Y sky130_fd_sc_hd__nor2_1
X_1947_ _1947_/A VGND VGND VPWR VPWR _2495_/A sky130_fd_sc_hd__inv_2
X_1878_ _1878_/A _1878_/B VGND VGND VPWR VPWR _1878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2850_ _2851_/A _2254_/Y _2262_/A _2820_/A _2849_/Y VGND VGND VPWR VPWR _2850_/X
+ sky130_fd_sc_hd__a221o_1
X_1801_ _1588_/Y _1642_/A _2265_/A _1783_/X VGND VGND VPWR VPWR _1802_/A sky130_fd_sc_hd__a31o_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _2794_/A _2781_/B VGND VGND VPWR VPWR _2781_/Y sky130_fd_sc_hd__nor2_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ _1763_/A _1732_/B _1747_/C VGND VGND VPWR VPWR _1736_/B sky130_fd_sc_hd__or3_4
XFILLER_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1663_ _2076_/A VGND VGND VPWR VPWR _2042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3402_ _3404_/CLK _3402_/D input1/X VGND VGND VPWR VPWR _3403_/D sky130_fd_sc_hd__dfrtp_1
X_1594_ _3389_/Q VGND VGND VPWR VPWR _2178_/A sky130_fd_sc_hd__clkbuf_2
X_3333_ _2312_/Y _2307_/Y _3340_/S VGND VGND VPWR VPWR _3333_/X sky130_fd_sc_hd__mux2_1
X_3264_ _3076_/Y _3074_/Y _3351_/S VGND VGND VPWR VPWR _3264_/X sky130_fd_sc_hd__mux2_2
X_2215_ _2215_/A _2286_/B VGND VGND VPWR VPWR _2597_/B sky130_fd_sc_hd__nor2_2
X_3195_ _2835_/Y _2831_/Y _3346_/S VGND VGND VPWR VPWR _3195_/X sky130_fd_sc_hd__mux2_2
X_2146_ _2148_/B VGND VGND VPWR VPWR _3039_/B sky130_fd_sc_hd__inv_2
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2077_ _2785_/A VGND VGND VPWR VPWR _2400_/B sky130_fd_sc_hd__inv_2
X_2979_ _3032_/A VGND VGND VPWR VPWR _2979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ _1974_/X _2989_/B _1963_/X _2756_/B _1999_/X VGND VGND VPWR VPWR _2000_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2902_ _3004_/A VGND VGND VPWR VPWR _3042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2833_ _2960_/A VGND VGND VPWR VPWR _2833_/X sky130_fd_sc_hd__clkbuf_2
X_2764_ _2004_/B _2761_/X _2992_/B _2753_/X _2763_/X VGND VGND VPWR VPWR _2764_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1715_ _3386_/Q _1847_/A _1744_/A VGND VGND VPWR VPWR _1945_/A sky130_fd_sc_hd__o21ai_2
X_2695_ _2929_/A _2581_/A _2328_/X _2434_/A VGND VGND VPWR VPWR _2695_/X sky130_fd_sc_hd__o22a_1
X_1646_ _1691_/A _1683_/A VGND VGND VPWR VPWR _2400_/A sky130_fd_sc_hd__or2_4
X_1577_ _2578_/B VGND VGND VPWR VPWR _2993_/A sky130_fd_sc_hd__clkbuf_2
X_3316_ _2144_/Y _2139_/Y _3381_/S VGND VGND VPWR VPWR _3316_/X sky130_fd_sc_hd__mux2_2
X_3247_ _3020_/Y _3018_/Y _3381_/S VGND VGND VPWR VPWR _3247_/X sky130_fd_sc_hd__mux2_1
X_3178_ _2771_/Y _2769_/Y _3370_/S VGND VGND VPWR VPWR _3178_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2129_ _2132_/B VGND VGND VPWR VPWR _3033_/B sky130_fd_sc_hd__inv_2
XFILLER_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput119 _3152_/X VGND VGND VPWR VPWR output_thermometer_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput108 _3241_/X VGND VGND VPWR VPWR output_thermometer_o[113] sky130_fd_sc_hd__clkbuf_2
X_2480_ _2726_/B _2459_/X _2479_/X VGND VGND VPWR VPWR _2480_/Y sky130_fd_sc_hd__o21ai_1
Xoutput90 _3300_/X VGND VGND VPWR VPWR output_thermometer_o[172] sky130_fd_sc_hd__clkbuf_2
X_3101_ _3101_/A VGND VGND VPWR VPWR _3101_/Y sky130_fd_sc_hd__inv_2
X_3032_ _3032_/A VGND VGND VPWR VPWR _3032_/X sky130_fd_sc_hd__buf_2
XFILLER_63_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2816_ _3022_/B VGND VGND VPWR VPWR _2854_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2747_ _2785_/C _2980_/B VGND VGND VPWR VPWR _2747_/X sky130_fd_sc_hd__or2_1
X_2678_ _2910_/B _2545_/X _2677_/X VGND VGND VPWR VPWR _2678_/Y sky130_fd_sc_hd__o21ai_1
X_1629_ _1683_/A VGND VGND VPWR VPWR _2044_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1980_ _1980_/A VGND VGND VPWR VPWR _2318_/A sky130_fd_sc_hd__clkinv_4
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2601_ _2766_/A VGND VGND VPWR VPWR _2723_/A sky130_fd_sc_hd__clkbuf_2
X_2532_ _2523_/X _3003_/B _3005_/B _2531_/X VGND VGND VPWR VPWR _2532_/X sky130_fd_sc_hd__o22a_1
X_2463_ _2949_/B VGND VGND VPWR VPWR _2463_/Y sky130_fd_sc_hd__inv_2
X_2394_ _1928_/A _2184_/A _2537_/A _2023_/X VGND VGND VPWR VPWR _3120_/A sky130_fd_sc_hd__a31o_1
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3015_ _3032_/A VGND VGND VPWR VPWR _3015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1963_ _2025_/A VGND VGND VPWR VPWR _1963_/X sky130_fd_sc_hd__clkbuf_2
X_1894_ _1854_/X _2955_/B _1842_/X _2722_/B _1893_/X VGND VGND VPWR VPWR _1894_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2515_ _2990_/B VGND VGND VPWR VPWR _2515_/Y sky130_fd_sc_hd__inv_2
X_2446_ _2446_/A _2785_/B VGND VGND VPWR VPWR _2936_/B sky130_fd_sc_hd__or2_2
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2377_ _2398_/A _2660_/A VGND VGND VPWR VPWR _3118_/B sky130_fd_sc_hd__or2_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3280_ _1676_/Y _1651_/Y _3347_/S VGND VGND VPWR VPWR _3280_/X sky130_fd_sc_hd__mux2_1
X_2300_ _3091_/B VGND VGND VPWR VPWR _2300_/Y sky130_fd_sc_hd__inv_2
X_2231_ _2400_/A _2231_/B VGND VGND VPWR VPWR _2236_/A sky130_fd_sc_hd__or2_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2162_ _2391_/C VGND VGND VPWR VPWR _2301_/C sky130_fd_sc_hd__buf_1
XFILLER_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2093_ _2093_/A _3022_/A VGND VGND VPWR VPWR _2096_/B sky130_fd_sc_hd__nand2_2
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2995_ _2978_/X _2004_/B _2979_/X _2760_/B _2994_/X VGND VGND VPWR VPWR _2995_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1946_ _1981_/A _2295_/A VGND VGND VPWR VPWR _1947_/A sky130_fd_sc_hd__or2_2
X_1877_ _1880_/B VGND VGND VPWR VPWR _1878_/B sky130_fd_sc_hd__inv_2
X_2429_ _2422_/X _2919_/B _2922_/A _2415_/X VGND VGND VPWR VPWR _2429_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1800_ _2178_/A VGND VGND VPWR VPWR _2265_/A sky130_fd_sc_hd__clkbuf_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _2867_/A VGND VGND VPWR VPWR _2794_/A sky130_fd_sc_hd__clkbuf_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ _2141_/B VGND VGND VPWR VPWR _1732_/B sky130_fd_sc_hd__inv_2
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1662_ _2178_/B VGND VGND VPWR VPWR _2076_/A sky130_fd_sc_hd__buf_2
X_3401_ _3404_/CLK _3401_/D input1/X VGND VGND VPWR VPWR _3402_/D sky130_fd_sc_hd__dfrtp_1
X_1593_ _1761_/A VGND VGND VPWR VPWR _2347_/A sky130_fd_sc_hd__clkbuf_2
X_3332_ _2305_/Y _2300_/Y _3340_/S VGND VGND VPWR VPWR _3332_/X sky130_fd_sc_hd__mux2_1
X_3263_ _3073_/Y _3071_/Y _3351_/S VGND VGND VPWR VPWR _3263_/X sky130_fd_sc_hd__mux2_2
X_3194_ _2830_/Y _2828_/Y _3346_/S VGND VGND VPWR VPWR _3194_/X sky130_fd_sc_hd__mux2_2
X_2214_ _2215_/A _2340_/A VGND VGND VPWR VPWR _3056_/B sky130_fd_sc_hd__nor2_2
X_2145_ _2042_/A _2310_/A _1684_/A _1605_/B VGND VGND VPWR VPWR _2148_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2076_ _2076_/A _2076_/B VGND VGND VPWR VPWR _2785_/A sky130_fd_sc_hd__nand2_2
XFILLER_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2978_ _3001_/A VGND VGND VPWR VPWR _2978_/X sky130_fd_sc_hd__clkbuf_2
X_1929_ _1978_/A _2486_/A _1954_/C VGND VGND VPWR VPWR _1929_/X sky130_fd_sc_hd__or3_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2901_ _2920_/A VGND VGND VPWR VPWR _2901_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2832_ _2832_/A VGND VGND VPWR VPWR _2960_/A sky130_fd_sc_hd__clkbuf_2
X_2763_ _2763_/A VGND VGND VPWR VPWR _2763_/X sky130_fd_sc_hd__clkbuf_2
X_1714_ _1581_/X _2681_/B _1713_/X VGND VGND VPWR VPWR _1714_/Y sky130_fd_sc_hd__o21ai_1
X_2694_ _2694_/A _2694_/B VGND VGND VPWR VPWR _2694_/Y sky130_fd_sc_hd__nor2_1
X_1645_ _2113_/A VGND VGND VPWR VPWR _1691_/A sky130_fd_sc_hd__inv_2
X_1576_ _2572_/A _3102_/A VGND VGND VPWR VPWR _2578_/B sky130_fd_sc_hd__or2_1
X_3315_ _2136_/Y _2130_/Y _3380_/S VGND VGND VPWR VPWR _3315_/X sky130_fd_sc_hd__mux2_1
X_3246_ _3017_/Y _3014_/Y _3374_/S VGND VGND VPWR VPWR _3246_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3177_ _2768_/Y _2765_/Y _3374_/S VGND VGND VPWR VPWR _3177_/X sky130_fd_sc_hd__mux2_2
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2128_ _2042_/A _2295_/A _1684_/A _1605_/B VGND VGND VPWR VPWR _2132_/B sky130_fd_sc_hd__a31o_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ _1992_/X _2019_/X _2020_/X _2534_/A _2023_/X VGND VGND VPWR VPWR _3008_/B
+ sky130_fd_sc_hd__o41a_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput109 _3201_/X VGND VGND VPWR VPWR output_thermometer_o[73] sky130_fd_sc_hd__clkbuf_2
Xoutput91 _3325_/X VGND VGND VPWR VPWR output_thermometer_o[197] sky130_fd_sc_hd__clkbuf_2
X_3100_ _3097_/X _2871_/B _3098_/X _2640_/B _3099_/X VGND VGND VPWR VPWR _3100_/Y
+ sky130_fd_sc_hd__o221ai_1
Xoutput80 _3249_/X VGND VGND VPWR VPWR output_thermometer_o[121] sky130_fd_sc_hd__clkbuf_2
X_3031_ _3041_/A _3031_/B VGND VGND VPWR VPWR _3031_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2815_ _2815_/A _2993_/A VGND VGND VPWR VPWR _3022_/B sky130_fd_sc_hd__or2_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2746_ _2756_/A _2746_/B VGND VGND VPWR VPWR _2746_/Y sky130_fd_sc_hd__nor2_1
X_2677_ _2911_/A _2611_/X _2393_/X _2413_/A VGND VGND VPWR VPWR _2677_/X sky130_fd_sc_hd__o22a_1
X_1628_ _1769_/B VGND VGND VPWR VPWR _1725_/B sky130_fd_sc_hd__clkbuf_2
X_3229_ _2954_/Y _2952_/Y _3357_/S VGND VGND VPWR VPWR _3229_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2600_ _2610_/A _2600_/B VGND VGND VPWR VPWR _2600_/Y sky130_fd_sc_hd__nor2_1
X_2531_ _2531_/A VGND VGND VPWR VPWR _2531_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2462_ _2462_/A _2471_/B VGND VGND VPWR VPWR _2949_/B sky130_fd_sc_hd__or2_2
X_2393_ _2785_/C VGND VGND VPWR VPWR _2393_/X sky130_fd_sc_hd__buf_2
XFILLER_68_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3014_ _3024_/A _3014_/B VGND VGND VPWR VPWR _3014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2729_ _1899_/B _2723_/X _2958_/B _2715_/X _2728_/X VGND VGND VPWR VPWR _2729_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ _1951_/X _2298_/B _1961_/X VGND VGND VPWR VPWR _2977_/B sky130_fd_sc_hd__a21oi_4
X_1893_ _1917_/A _2471_/A _1893_/C VGND VGND VPWR VPWR _1893_/X sky130_fd_sc_hd__or3_2
X_2514_ _2514_/A _2514_/B VGND VGND VPWR VPWR _2990_/B sky130_fd_sc_hd__or2_2
X_2445_ _2324_/X _1799_/Y _2444_/X VGND VGND VPWR VPWR _2445_/Y sky130_fd_sc_hd__o21ai_1
X_2376_ _2103_/A _2058_/A _2009_/B VGND VGND VPWR VPWR _2660_/A sky130_fd_sc_hd__o21a_1
XFILLER_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput270 _3363_/X VGND VGND VPWR VPWR output_thermometer_o[235] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2230_ _3065_/B VGND VGND VPWR VPWR _2230_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2161_ _2161_/A VGND VGND VPWR VPWR _2161_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2092_ _2103_/A _2548_/A _2092_/C VGND VGND VPWR VPWR _3022_/A sky130_fd_sc_hd__or3_4
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2994_ _2994_/A VGND VGND VPWR VPWR _2994_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1945_ _1945_/A VGND VGND VPWR VPWR _2295_/A sky130_fd_sc_hd__inv_4
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1876_ _1871_/X _2467_/A _1875_/X VGND VGND VPWR VPWR _1880_/B sky130_fd_sc_hd__o21ai_2
X_2428_ _2527_/A VGND VGND VPWR VPWR _2428_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2359_ _2359_/A _2654_/A VGND VGND VPWR VPWR _3112_/B sky130_fd_sc_hd__or2_2
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1730_ _1884_/A _1759_/A _1761_/A VGND VGND VPWR VPWR _2141_/B sky130_fd_sc_hd__or3_4
X_1661_ _1661_/A VGND VGND VPWR VPWR _2178_/B sky130_fd_sc_hd__inv_2
X_3400_ _3404_/CLK _3400_/D input1/X VGND VGND VPWR VPWR _3401_/D sky130_fd_sc_hd__dfrtp_1
X_1592_ _1661_/A VGND VGND VPWR VPWR _1761_/A sky130_fd_sc_hd__buf_1
X_3331_ _2297_/Y _2290_/Y _3340_/S VGND VGND VPWR VPWR _3331_/X sky130_fd_sc_hd__mux2_1
X_3262_ _3070_/Y _3068_/Y _3330_/S VGND VGND VPWR VPWR _3262_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2213_ _2184_/X _3058_/B _2185_/X VGND VGND VPWR VPWR _2831_/B sky130_fd_sc_hd__o21a_1
X_3193_ _2827_/Y _2823_/Y _3330_/S VGND VGND VPWR VPWR _3193_/X sky130_fd_sc_hd__mux2_2
X_2144_ _2131_/X _2805_/B _2143_/X VGND VGND VPWR VPWR _2144_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2075_ _2109_/A _2075_/B VGND VGND VPWR VPWR _2075_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2977_ _2985_/A _2977_/B VGND VGND VPWR VPWR _2977_/Y sky130_fd_sc_hd__nor2_1
X_1928_ _1928_/A VGND VGND VPWR VPWR _1978_/A sky130_fd_sc_hd__clkbuf_2
X_1859_ _1854_/X _2945_/B _1842_/X _2711_/B _1858_/X VGND VGND VPWR VPWR _1859_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_1_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2900_ _2905_/A _2900_/B VGND VGND VPWR VPWR _2900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2831_ _2839_/A _2831_/B VGND VGND VPWR VPWR _2831_/Y sky130_fd_sc_hd__nor2_1
X_2762_ _2762_/A _2993_/B VGND VGND VPWR VPWR _2763_/A sky130_fd_sc_hd__or2_1
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ _1708_/X _2418_/A _1622_/X _2913_/B VGND VGND VPWR VPWR _1713_/X sky130_fd_sc_hd__o22a_1
XANTENNA_0 _2948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2693_ _2924_/B _2682_/X _2692_/X VGND VGND VPWR VPWR _2693_/Y sky130_fd_sc_hd__o21ai_1
X_1644_ _1884_/A VGND VGND VPWR VPWR _2548_/A sky130_fd_sc_hd__buf_2
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1575_ input2/X _3408_/Q VGND VGND VPWR VPWR _3102_/A sky130_fd_sc_hd__nand2_2
X_3314_ _2127_/Y _2121_/Y _3380_/S VGND VGND VPWR VPWR _3314_/X sky130_fd_sc_hd__mux2_1
X_3245_ _3013_/Y _3011_/Y _3381_/S VGND VGND VPWR VPWR _3245_/X sky130_fd_sc_hd__mux2_1
X_3176_ _2764_/Y _2760_/Y _3370_/S VGND VGND VPWR VPWR _3176_/X sky130_fd_sc_hd__mux2_2
X_2127_ _1735_/X _2798_/B _2126_/X VGND VGND VPWR VPWR _2127_/Y sky130_fd_sc_hd__o21ai_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ _2058_/A VGND VGND VPWR VPWR _2534_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput70 _3373_/X VGND VGND VPWR VPWR output_thermometer_o[245] sky130_fd_sc_hd__clkbuf_2
Xoutput81 _3314_/X VGND VGND VPWR VPWR output_thermometer_o[186] sky130_fd_sc_hd__clkbuf_2
Xoutput92 _3360_/X VGND VGND VPWR VPWR output_thermometer_o[232] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3030_ _2800_/A _2920_/X _3015_/X _2798_/B _3029_/X VGND VGND VPWR VPWR _3030_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2814_ _2165_/B _2577_/A _3044_/A _2577_/B VGND VGND VPWR VPWR _2814_/X sky130_fd_sc_hd__o211a_1
X_2745_ _1950_/B _2743_/X _2974_/B _2734_/X _2744_/X VGND VGND VPWR VPWR _2745_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2676_ _2676_/A _2676_/B VGND VGND VPWR VPWR _2676_/Y sky130_fd_sc_hd__nor2_1
X_1627_ _1627_/A VGND VGND VPWR VPWR _1769_/B sky130_fd_sc_hd__buf_2
X_3228_ _2950_/Y _2948_/Y _3357_/S VGND VGND VPWR VPWR _3228_/X sky130_fd_sc_hd__mux2_1
X_3159_ _2699_/Y _2697_/Y _3351_/S VGND VGND VPWR VPWR _3159_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _2530_/A _2548_/B VGND VGND VPWR VPWR _2530_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2461_ _2711_/B _2459_/X _2460_/X VGND VGND VPWR VPWR _2461_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2392_ _2762_/A VGND VGND VPWR VPWR _2785_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3013_ _1797_/X _2538_/A _2997_/X _2781_/B _3012_/X VGND VGND VPWR VPWR _3013_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2728_ _2744_/A _2962_/B VGND VGND VPWR VPWR _2728_/X sky130_fd_sc_hd__or2_1
X_2659_ _2659_/A _2659_/B VGND VGND VPWR VPWR _2659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1961_ _2193_/A VGND VGND VPWR VPWR _1961_/X sky130_fd_sc_hd__buf_4
X_1892_ _1903_/A _1892_/B VGND VGND VPWR VPWR _2722_/B sky130_fd_sc_hd__nor2_2
X_2513_ _2752_/B _2506_/X _2512_/X VGND VGND VPWR VPWR _2513_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2444_ _2341_/X _1794_/Y _2301_/A _2436_/X VGND VGND VPWR VPWR _2444_/X sky130_fd_sc_hd__o22a_1
X_2375_ _2351_/X _2656_/B _2374_/X VGND VGND VPWR VPWR _2375_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput260 _3208_/X VGND VGND VPWR VPWR output_thermometer_o[80] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2160_ _2131_/X _2811_/B _2159_/X VGND VGND VPWR VPWR _2160_/Y sky130_fd_sc_hd__o21ai_1
X_2091_ _2087_/X _3018_/B _2080_/X _2787_/B _2090_/X VGND VGND VPWR VPWR _2091_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2993_ _2993_/A _2993_/B VGND VGND VPWR VPWR _2994_/A sky130_fd_sc_hd__or2_1
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1944_ _3047_/A VGND VGND VPWR VPWR _1996_/A sky130_fd_sc_hd__clkbuf_2
X_1875_ _2233_/A VGND VGND VPWR VPWR _1875_/X sky130_fd_sc_hd__buf_2
X_2427_ _2791_/A VGND VGND VPWR VPWR _2527_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2358_ _2347_/X _2036_/A _2009_/B VGND VGND VPWR VPWR _2654_/A sky130_fd_sc_hd__o21a_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2289_ _2295_/A _2289_/B VGND VGND VPWR VPWR _3088_/B sky130_fd_sc_hd__nor2_2
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1660_ _3097_/A VGND VGND VPWR VPWR _1660_/X sky130_fd_sc_hd__buf_2
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1591_ _1588_/Y _1570_/A _1991_/A VGND VGND VPWR VPWR _1661_/A sky130_fd_sc_hd__o21ai_1
X_3330_ _2288_/Y _2283_/Y _3330_/S VGND VGND VPWR VPWR _3330_/X sky130_fd_sc_hd__mux2_2
X_3261_ _3066_/Y _3064_/Y _3330_/S VGND VGND VPWR VPWR _3261_/X sky130_fd_sc_hd__mux2_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3192_ _2821_/Y _1792_/A _3346_/S VGND VGND VPWR VPWR _3192_/X sky130_fd_sc_hd__mux2_2
X_2212_ _2315_/A VGND VGND VPWR VPWR _2212_/X sky130_fd_sc_hd__clkbuf_2
X_2143_ _1818_/A _3035_/B _2141_/B _1802_/X VGND VGND VPWR VPWR _2143_/X sky130_fd_sc_hd__o22a_1
X_2074_ _2081_/B VGND VGND VPWR VPWR _2075_/B sky130_fd_sc_hd__inv_2
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2976_ _2959_/X _1950_/B _2960_/X _2741_/B _2975_/X VGND VGND VPWR VPWR _2976_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1927_ _1964_/A _1927_/B VGND VGND VPWR VPWR _2733_/B sky130_fd_sc_hd__nor2_4
X_1858_ _1858_/A _2457_/A _1893_/C VGND VGND VPWR VPWR _1858_/X sky130_fd_sc_hd__or3_2
X_1789_ _2705_/A VGND VGND VPWR VPWR _1789_/X sky130_fd_sc_hd__buf_2
XFILLER_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2830_ _2825_/X _3051_/B _1660_/X _2593_/B _2829_/X VGND VGND VPWR VPWR _2830_/Y
+ sky130_fd_sc_hd__o221ai_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ _2920_/A VGND VGND VPWR VPWR _2761_/X sky130_fd_sc_hd__clkbuf_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2692_ _2925_/A _2581_/A _2328_/X _2431_/A VGND VGND VPWR VPWR _2692_/X sky130_fd_sc_hd__o22a_1
X_1712_ _1725_/A _1725_/B _1712_/C VGND VGND VPWR VPWR _2913_/B sky130_fd_sc_hd__and3_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1643_ _1664_/A VGND VGND VPWR VPWR _1884_/A sky130_fd_sc_hd__inv_2
XANTENNA_1 _3377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ _1618_/A VGND VGND VPWR VPWR _2572_/A sky130_fd_sc_hd__inv_2
X_3313_ _2117_/Y _2109_/Y _3381_/S VGND VGND VPWR VPWR _3313_/X sky130_fd_sc_hd__mux2_1
X_3244_ _3010_/Y _3008_/Y _3370_/S VGND VGND VPWR VPWR _3244_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3175_ _2758_/Y _2756_/Y _3370_/S VGND VGND VPWR VPWR _3175_/X sky130_fd_sc_hd__mux2_2
X_2126_ _1755_/X _3028_/B _2124_/B _1802_/X VGND VGND VPWR VPWR _2126_/X sky130_fd_sc_hd__o22a_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2057_ _2057_/A VGND VGND VPWR VPWR _2058_/A sky130_fd_sc_hd__inv_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2959_ _3001_/A VGND VGND VPWR VPWR _2959_/X sky130_fd_sc_hd__buf_2
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput60 _3343_/X VGND VGND VPWR VPWR output_thermometer_o[215] sky130_fd_sc_hd__clkbuf_2
Xoutput71 _3210_/X VGND VGND VPWR VPWR output_thermometer_o[82] sky130_fd_sc_hd__clkbuf_2
Xoutput93 _3370_/X VGND VGND VPWR VPWR output_thermometer_o[242] sky130_fd_sc_hd__clkbuf_2
Xoutput82 _3340_/X VGND VGND VPWR VPWR output_thermometer_o[212] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2813_ _3042_/B _2799_/X _3041_/B _2256_/X _2812_/X VGND VGND VPWR VPWR _2813_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_8_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2744_ _2744_/A _2975_/B VGND VGND VPWR VPWR _2744_/X sky130_fd_sc_hd__or2_1
X_2675_ _2907_/A _2653_/X _2905_/B _2673_/X _2674_/X VGND VGND VPWR VPWR _2675_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1626_ _1722_/A VGND VGND VPWR VPWR _1725_/A sky130_fd_sc_hd__clkbuf_2
X_3227_ _2947_/Y _2945_/Y _3354_/S VGND VGND VPWR VPWR _3227_/X sky130_fd_sc_hd__mux2_4
X_3158_ _2696_/Y _2694_/Y _3380_/S VGND VGND VPWR VPWR _3158_/X sky130_fd_sc_hd__mux2_1
X_2109_ _2109_/A _3025_/B VGND VGND VPWR VPWR _2109_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3089_ _3078_/X _2861_/B _3079_/X _2629_/B _3088_/X VGND VGND VPWR VPWR _3089_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2460_ _2454_/X _2945_/B _1852_/B _2436_/X VGND VGND VPWR VPWR _2460_/X sky130_fd_sc_hd__o22a_1
X_2391_ _2391_/A _2537_/A _2391_/C VGND VGND VPWR VPWR _2663_/B sky130_fd_sc_hd__and3_1
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3012_ _3029_/A _3012_/B VGND VGND VPWR VPWR _3012_/X sky130_fd_sc_hd__or2_1
X_2727_ _2727_/A VGND VGND VPWR VPWR _2744_/A sky130_fd_sc_hd__buf_1
X_2658_ _3114_/B _2653_/X _2171_/A _2886_/B _2657_/X VGND VGND VPWR VPWR _2658_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2589_ _2589_/A VGND VGND VPWR VPWR _2618_/B sky130_fd_sc_hd__clkbuf_2
X_1609_ _3057_/A VGND VGND VPWR VPWR _3099_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1960_ _1996_/A _1960_/B VGND VGND VPWR VPWR _1960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1891_ _1890_/X _2243_/B _1840_/X VGND VGND VPWR VPWR _2955_/B sky130_fd_sc_hd__a21oi_4
X_2512_ _2501_/X _2985_/B _1985_/B _2511_/X VGND VGND VPWR VPWR _2512_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2443_ _2785_/B VGND VGND VPWR VPWR _2443_/Y sky130_fd_sc_hd__inv_2
X_2374_ _2246_/X _2886_/B _2248_/X _3114_/B VGND VGND VPWR VPWR _2374_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput261 _3135_/X VGND VGND VPWR VPWR output_thermometer_o[7] sky130_fd_sc_hd__clkbuf_2
Xoutput250 _3250_/X VGND VGND VPWR VPWR output_thermometer_o[122] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2090_ _2090_/A _2090_/B VGND VGND VPWR VPWR _2090_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2992_ _3003_/A _2992_/B VGND VGND VPWR VPWR _2992_/Y sky130_fd_sc_hd__nor2_1
X_1943_ _2898_/A VGND VGND VPWR VPWR _3047_/A sky130_fd_sc_hd__clkbuf_4
X_1874_ _2231_/B VGND VGND VPWR VPWR _2467_/A sky130_fd_sc_hd__inv_2
X_2426_ _2426_/A VGND VGND VPWR VPWR _2791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2357_ _2351_/X _2649_/B _2356_/X VGND VGND VPWR VPWR _2357_/Y sky130_fd_sc_hd__o21ai_1
X_2288_ _2212_/X _2856_/B _2287_/X VGND VGND VPWR VPWR _2288_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ _1860_/A _1642_/A VGND VGND VPWR VPWR _1991_/A sky130_fd_sc_hd__or2_2
X_3260_ _3063_/Y _3060_/Y _3346_/S VGND VGND VPWR VPWR _3260_/X sky130_fd_sc_hd__mux2_2
X_3191_ _2814_/X _2166_/X _3365_/S VGND VGND VPWR VPWR _3191_/X sky130_fd_sc_hd__mux2_2
X_2211_ _2290_/A _3058_/B VGND VGND VPWR VPWR _2211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2142_ _2142_/A _2806_/A VGND VGND VPWR VPWR _3035_/B sky130_fd_sc_hd__and2_1
X_2073_ _2005_/X _2076_/B _2397_/A _2014_/X VGND VGND VPWR VPWR _2081_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2975_ _2975_/A _2975_/B VGND VGND VPWR VPWR _2975_/X sky130_fd_sc_hd__or2_1
X_1926_ _1890_/X _1922_/A _1900_/X VGND VGND VPWR VPWR _2967_/B sky130_fd_sc_hd__a21oi_4
X_1857_ _1903_/A _1857_/B VGND VGND VPWR VPWR _2711_/B sky130_fd_sc_hd__nor2_4
X_1788_ _2727_/A VGND VGND VPWR VPWR _2705_/A sky130_fd_sc_hd__clkbuf_2
X_2409_ _2669_/B _2171_/X _2408_/X VGND VGND VPWR VPWR _2409_/Y sky130_fd_sc_hd__o21ai_1
X_3389_ _3408_/CLK _3389_/D VGND VGND VPWR VPWR _3389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ _2776_/A _2760_/B VGND VGND VPWR VPWR _2760_/Y sky130_fd_sc_hd__nor2_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2691_ _2694_/A _2691_/B VGND VGND VPWR VPWR _2691_/Y sky130_fd_sc_hd__nor2_1
X_1711_ _1769_/A _1712_/C VGND VGND VPWR VPWR _2418_/A sky130_fd_sc_hd__or2_2
XANTENNA_2 _3207_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _1642_/A _2617_/A VGND VGND VPWR VPWR _1664_/A sky130_fd_sc_hd__or2_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1573_ input2/X _3408_/D VGND VGND VPWR VPWR _1618_/A sky130_fd_sc_hd__nand2_1
X_3312_ _2106_/Y _2095_/Y _3381_/S VGND VGND VPWR VPWR _3312_/X sky130_fd_sc_hd__mux2_1
X_3243_ _3006_/Y _3003_/Y _3370_/S VGND VGND VPWR VPWR _3243_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3174_ _2755_/Y _2752_/Y _3370_/S VGND VGND VPWR VPWR _3174_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2125_ _2158_/A _2800_/A VGND VGND VPWR VPWR _3028_/B sky130_fd_sc_hd__and2_1
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2056_ _2056_/A _3009_/B VGND VGND VPWR VPWR _2056_/Y sky130_fd_sc_hd__nor2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2958_ _2967_/A _2958_/B VGND VGND VPWR VPWR _2958_/Y sky130_fd_sc_hd__nor2_1
X_1909_ _1909_/A VGND VGND VPWR VPWR _2481_/A sky130_fd_sc_hd__inv_2
X_2889_ _2889_/A VGND VGND VPWR VPWR _2970_/A sky130_fd_sc_hd__buf_2
XFILLER_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput50 _3230_/X VGND VGND VPWR VPWR output_thermometer_o[102] sky130_fd_sc_hd__clkbuf_2
Xoutput61 _3220_/X VGND VGND VPWR VPWR output_thermometer_o[92] sky130_fd_sc_hd__clkbuf_2
Xoutput72 _3308_/X VGND VGND VPWR VPWR output_thermometer_o[180] sky130_fd_sc_hd__clkbuf_2
Xoutput83 _3322_/X VGND VGND VPWR VPWR output_thermometer_o[194] sky130_fd_sc_hd__clkbuf_2
Xoutput94 _3331_/X VGND VGND VPWR VPWR output_thermometer_o[203] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2812_ _2812_/A _2849_/A VGND VGND VPWR VPWR _2812_/X sky130_fd_sc_hd__or2_1
X_2743_ _2920_/A VGND VGND VPWR VPWR _2743_/X sky130_fd_sc_hd__clkbuf_2
X_2674_ _2674_/A _2803_/B VGND VGND VPWR VPWR _2674_/X sky130_fd_sc_hd__or2_1
X_1625_ _2578_/A VGND VGND VPWR VPWR _1722_/A sky130_fd_sc_hd__clkbuf_2
X_3226_ _2944_/Y _2938_/Y _3354_/S VGND VGND VPWR VPWR _3226_/X sky130_fd_sc_hd__mux2_1
X_3157_ _2693_/Y _2691_/Y _3347_/S VGND VGND VPWR VPWR _3157_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2108_ _2111_/B VGND VGND VPWR VPWR _3025_/B sky130_fd_sc_hd__inv_2
XFILLER_54_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3088_ _3099_/A _3088_/B _3094_/C VGND VGND VPWR VPWR _3088_/X sky130_fd_sc_hd__or3_1
X_2039_ _2081_/A _2039_/B VGND VGND VPWR VPWR _2769_/B sky130_fd_sc_hd__nor2_2
XFILLER_22_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2390_ _2390_/A VGND VGND VPWR VPWR _2390_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3011_ _3024_/A _3011_/B VGND VGND VPWR VPWR _3011_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2726_ _2737_/A _2726_/B VGND VGND VPWR VPWR _2726_/Y sky130_fd_sc_hd__nor2_1
X_2657_ _2657_/A _2660_/B VGND VGND VPWR VPWR _2657_/X sky130_fd_sc_hd__or2_1
X_1608_ _2168_/A VGND VGND VPWR VPWR _3057_/A sky130_fd_sc_hd__buf_1
X_2588_ _2931_/A _2588_/B VGND VGND VPWR VPWR _2588_/Y sky130_fd_sc_hd__nor2_1
X_3209_ _2880_/Y _2878_/Y _3340_/S VGND VGND VPWR VPWR _3209_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1890_ _1890_/A VGND VGND VPWR VPWR _1890_/X sky130_fd_sc_hd__buf_4
X_2511_ _2531_/A VGND VGND VPWR VPWR _2511_/X sky130_fd_sc_hd__clkbuf_2
X_2442_ _2514_/B VGND VGND VPWR VPWR _2785_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2373_ _2373_/A VGND VGND VPWR VPWR _3114_/B sky130_fd_sc_hd__inv_2
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2709_ _2724_/A _2943_/B VGND VGND VPWR VPWR _2709_/X sky130_fd_sc_hd__or2_1
Xoutput251 _3129_/X VGND VGND VPWR VPWR output_thermometer_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput240 _3184_/X VGND VGND VPWR VPWR output_thermometer_o[56] sky130_fd_sc_hd__clkbuf_2
Xoutput262 _3203_/X VGND VGND VPWR VPWR output_thermometer_o[75] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2991_ _2978_/X _1996_/B _2979_/X _2756_/B _2990_/X VGND VGND VPWR VPWR _2991_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1942_ _1913_/X _2971_/B _1902_/X _2737_/B _1941_/X VGND VGND VPWR VPWR _1942_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_61_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1873_ _1907_/A _2067_/B VGND VGND VPWR VPWR _2231_/B sky130_fd_sc_hd__or2_4
X_2425_ _2425_/A VGND VGND VPWR VPWR _2425_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2356_ _2246_/X _2878_/B _2248_/X _3107_/B VGND VGND VPWR VPWR _2356_/X sky130_fd_sc_hd__o22a_1
X_2287_ _2263_/A _3083_/B _2606_/A _2625_/B VGND VGND VPWR VPWR _2287_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2210_ _2215_/A _2289_/B VGND VGND VPWR VPWR _3058_/B sky130_fd_sc_hd__nor2_2
X_3190_ _2813_/Y _2811_/Y _3382_/S VGND VGND VPWR VPWR _3190_/X sky130_fd_sc_hd__mux2_2
X_2141_ _2149_/A _2141_/B _2141_/C VGND VGND VPWR VPWR _2806_/A sky130_fd_sc_hd__or3_4
X_2072_ _2034_/X _3011_/B _2025_/X _2781_/B _2071_/X VGND VGND VPWR VPWR _2072_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2974_ _2985_/A _2974_/B VGND VGND VPWR VPWR _2974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1925_ _1938_/A _1925_/B VGND VGND VPWR VPWR _1925_/Y sky130_fd_sc_hd__nor2_1
X_1856_ _2038_/A VGND VGND VPWR VPWR _1903_/A sky130_fd_sc_hd__buf_4
X_1787_ _2762_/A VGND VGND VPWR VPWR _2727_/A sky130_fd_sc_hd__clkbuf_2
X_2408_ _2381_/X _2900_/B _3126_/B _2173_/X VGND VGND VPWR VPWR _2408_/X sky130_fd_sc_hd__o22a_1
X_3388_ _3408_/CLK input9/X VGND VGND VPWR VPWR _3388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2339_ _3080_/A _3105_/B VGND VGND VPWR VPWR _2339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ _2919_/B _2682_/X _2689_/X VGND VGND VPWR VPWR _2690_/Y sky130_fd_sc_hd__o21ai_1
X_1710_ _2386_/A _1704_/B _1709_/X VGND VGND VPWR VPWR _1712_/C sky130_fd_sc_hd__o21ai_1
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _3373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1641_ _2788_/A _1641_/B VGND VGND VPWR VPWR _2617_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3311_ _2091_/Y _2086_/Y _3381_/S VGND VGND VPWR VPWR _3311_/X sky130_fd_sc_hd__mux2_1
X_1572_ _1627_/A VGND VGND VPWR VPWR _2168_/B sky130_fd_sc_hd__inv_2
X_3242_ _3002_/Y _3000_/Y _3370_/S VGND VGND VPWR VPWR _3242_/X sky130_fd_sc_hd__mux2_1
X_3173_ _2751_/Y _2749_/Y _3370_/S VGND VGND VPWR VPWR _3173_/X sky130_fd_sc_hd__mux2_2
X_2124_ _2149_/A _2124_/B _2141_/C VGND VGND VPWR VPWR _2800_/A sky130_fd_sc_hd__or3_4
XFILLER_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2055_ _2060_/B VGND VGND VPWR VPWR _3009_/B sky130_fd_sc_hd__inv_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2957_ _2940_/X _1889_/B _2941_/X _2722_/B _2956_/X VGND VGND VPWR VPWR _2957_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1908_ _2265_/B _2268_/B VGND VGND VPWR VPWR _1909_/A sky130_fd_sc_hd__or2_4
X_2888_ _2882_/X _2656_/B _2840_/X _3115_/B _2887_/X VGND VGND VPWR VPWR _2888_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1839_ _1839_/A VGND VGND VPWR VPWR _1900_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput51 _3252_/X VGND VGND VPWR VPWR output_thermometer_o[124] sky130_fd_sc_hd__clkbuf_2
Xoutput40 _3206_/X VGND VGND VPWR VPWR output_thermometer_o[78] sky130_fd_sc_hd__clkbuf_2
Xoutput84 _3372_/X VGND VGND VPWR VPWR output_thermometer_o[244] sky130_fd_sc_hd__clkbuf_2
Xoutput73 _3182_/X VGND VGND VPWR VPWR output_thermometer_o[54] sky130_fd_sc_hd__clkbuf_2
Xoutput62 _3299_/X VGND VGND VPWR VPWR output_thermometer_o[171] sky130_fd_sc_hd__clkbuf_2
Xoutput95 _3223_/X VGND VGND VPWR VPWR output_thermometer_o[95] sky130_fd_sc_hd__clkbuf_2
XFILLER_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2811_ _2811_/A _2811_/B VGND VGND VPWR VPWR _2811_/Y sky130_fd_sc_hd__nor2_1
X_2742_ _2766_/A VGND VGND VPWR VPWR _2920_/A sky130_fd_sc_hd__buf_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2673_ _2715_/A VGND VGND VPWR VPWR _2673_/X sky130_fd_sc_hd__buf_2
X_1624_ _2391_/C _1624_/B VGND VGND VPWR VPWR _2578_/A sky130_fd_sc_hd__or2_2
X_3225_ _2937_/Y _2935_/Y _3351_/S VGND VGND VPWR VPWR _3225_/X sky130_fd_sc_hd__mux2_2
X_3156_ _2690_/Y _2688_/Y _3380_/S VGND VGND VPWR VPWR _3156_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2107_ _2042_/X _2279_/A _2030_/X _2044_/X VGND VGND VPWR VPWR _2111_/B sky130_fd_sc_hd__a31o_1
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3087_ _3107_/A _3087_/B VGND VGND VPWR VPWR _3087_/Y sky130_fd_sc_hd__nor2_1
X_2038_ _2038_/A VGND VGND VPWR VPWR _2081_/A sky130_fd_sc_hd__buf_4
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3010_ _2534_/A _2994_/X _2997_/X _2776_/B _3009_/X VGND VGND VPWR VPWR _3010_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_51_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2725_ _1889_/B _2723_/X _2955_/B _2715_/X _2724_/X VGND VGND VPWR VPWR _2725_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2656_ _2659_/A _2656_/B VGND VGND VPWR VPWR _2656_/Y sky130_fd_sc_hd__nor2_1
X_1607_ _1618_/A _3102_/A VGND VGND VPWR VPWR _2168_/A sky130_fd_sc_hd__or2_4
X_2587_ _2662_/A VGND VGND VPWR VPWR _2931_/A sky130_fd_sc_hd__buf_2
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3208_ _2877_/X _2343_/A _3354_/S VGND VGND VPWR VPWR _3208_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3139_ _2632_/Y _2629_/Y _3340_/S VGND VGND VPWR VPWR _3139_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2510_ _2986_/B VGND VGND VPWR VPWR _2510_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2441_ _2697_/B _2256_/X _2080_/X _2931_/B _2440_/X VGND VGND VPWR VPWR _2441_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2372_ _2233_/X _2657_/A _2234_/X VGND VGND VPWR VPWR _2886_/B sky130_fd_sc_hd__o21a_1
XFILLER_68_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2708_ _2727_/A VGND VGND VPWR VPWR _2724_/A sky130_fd_sc_hd__clkbuf_2
Xoutput241 _3247_/X VGND VGND VPWR VPWR output_thermometer_o[119] sky130_fd_sc_hd__clkbuf_2
X_2639_ _2662_/A VGND VGND VPWR VPWR _2659_/A sky130_fd_sc_hd__clkbuf_2
Xoutput252 _3279_/X VGND VGND VPWR VPWR output_thermometer_o[151] sky130_fd_sc_hd__clkbuf_2
Xoutput230 _3293_/X VGND VGND VPWR VPWR output_thermometer_o[165] sky130_fd_sc_hd__clkbuf_2
Xoutput263 _3375_/X VGND VGND VPWR VPWR output_thermometer_o[247] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2990_ _2990_/A _2990_/B VGND VGND VPWR VPWR _2990_/X sky130_fd_sc_hd__or2_1
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1941_ _1978_/A _2491_/A _1954_/C VGND VGND VPWR VPWR _1941_/X sky130_fd_sc_hd__or3_1
X_1872_ _2268_/B _1872_/B VGND VGND VPWR VPWR _2067_/B sky130_fd_sc_hd__or2_2
X_2424_ _2685_/B _2171_/X _2423_/X VGND VGND VPWR VPWR _2424_/Y sky130_fd_sc_hd__o21ai_1
X_2355_ _2355_/A VGND VGND VPWR VPWR _3107_/B sky130_fd_sc_hd__inv_2
X_2286_ _2286_/A _2286_/B VGND VGND VPWR VPWR _2625_/B sky130_fd_sc_hd__nor2_2
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2232_/A _2140_/B VGND VGND VPWR VPWR _2805_/B sky130_fd_sc_hd__nor2_4
X_2071_ _2082_/A _2537_/A _2071_/C VGND VGND VPWR VPWR _2071_/X sky130_fd_sc_hd__or3_1
XFILLER_61_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2973_ _2959_/X _1938_/B _2960_/X _2737_/B _2972_/X VGND VGND VPWR VPWR _2973_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1924_ _1927_/B VGND VGND VPWR VPWR _1925_/B sky130_fd_sc_hd__inv_2
X_1855_ _1820_/X _1849_/A _1840_/X VGND VGND VPWR VPWR _2945_/B sky130_fd_sc_hd__a21oi_4
X_1786_ _1786_/A _2301_/A VGND VGND VPWR VPWR _1786_/Y sky130_fd_sc_hd__nor2_1
X_2407_ _2407_/A VGND VGND VPWR VPWR _3126_/B sky130_fd_sc_hd__inv_2
X_3387_ _3408_/CLK input8/X VGND VGND VPWR VPWR _3387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2338_ _2338_/A VGND VGND VPWR VPWR _3105_/B sky130_fd_sc_hd__inv_2
X_2269_ _2269_/A VGND VGND VPWR VPWR _3074_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1640_ _3387_/Q VGND VGND VPWR VPWR _2788_/A sky130_fd_sc_hd__inv_2
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 _3213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1571_ _3391_/Q _1601_/A VGND VGND VPWR VPWR _1627_/A sky130_fd_sc_hd__or2_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3310_ _2083_/Y _2075_/Y _3381_/S VGND VGND VPWR VPWR _3310_/X sky130_fd_sc_hd__mux2_1
X_3241_ _2999_/Y _2996_/Y _3374_/S VGND VGND VPWR VPWR _3241_/X sky130_fd_sc_hd__mux2_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3172_ _2748_/Y _2746_/Y _3365_/S VGND VGND VPWR VPWR _3172_/X sky130_fd_sc_hd__mux2_2
X_2123_ _2234_/A VGND VGND VPWR VPWR _2158_/A sky130_fd_sc_hd__buf_1
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2054_ _2042_/X _2057_/A _2030_/X _2044_/X VGND VGND VPWR VPWR _2060_/B sky130_fd_sc_hd__a31o_1
XFILLER_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2956_ _2956_/A _2956_/B VGND VGND VPWR VPWR _2956_/X sky130_fd_sc_hd__or2_1
X_1907_ _1907_/A VGND VGND VPWR VPWR _2265_/B sky130_fd_sc_hd__clkbuf_2
X_2887_ _2887_/A _3114_/B _3049_/C VGND VGND VPWR VPWR _2887_/X sky130_fd_sc_hd__or3_2
X_1838_ _1878_/A _1838_/B VGND VGND VPWR VPWR _1838_/Y sky130_fd_sc_hd__nor2_1
X_1769_ _1769_/A _1769_/B _1769_/C VGND VGND VPWR VPWR _2928_/B sky130_fd_sc_hd__and3_1
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput41 _3244_/X VGND VGND VPWR VPWR output_thermometer_o[116] sky130_fd_sc_hd__clkbuf_2
Xoutput52 _3234_/X VGND VGND VPWR VPWR output_thermometer_o[106] sky130_fd_sc_hd__clkbuf_2
Xoutput30 _3200_/X VGND VGND VPWR VPWR output_thermometer_o[72] sky130_fd_sc_hd__clkbuf_2
Xoutput85 _3310_/X VGND VGND VPWR VPWR output_thermometer_o[182] sky130_fd_sc_hd__clkbuf_2
Xoutput63 _3222_/X VGND VGND VPWR VPWR output_thermometer_o[94] sky130_fd_sc_hd__clkbuf_2
Xoutput74 _3251_/X VGND VGND VPWR VPWR output_thermometer_o[123] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput96 _3258_/X VGND VGND VPWR VPWR output_thermometer_o[130] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2810_ _3039_/B _2799_/X _3038_/B _2256_/X _2809_/X VGND VGND VPWR VPWR _2810_/Y
+ sky130_fd_sc_hd__o221ai_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _2756_/A _2741_/B VGND VGND VPWR VPWR _2741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2672_ _2676_/A _2672_/B VGND VGND VPWR VPWR _2672_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1623_ _3391_/Q VGND VGND VPWR VPWR _2391_/C sky130_fd_sc_hd__inv_2
X_3224_ _2934_/Y _1794_/A _3342_/S VGND VGND VPWR VPWR _3224_/X sky130_fd_sc_hd__mux2_2
.ends

