**.subckt bandgap_core_test
**.ends
.end
