**.subckt bandgap_core_verification
xdut vdd ptat ctat cas GND en ctl_ptat[4] ctl_ptat[3] ctl_ptat[2] ctl_ptat[1] ctl_ptat[0]
+ ctl_ctat[4] ctl_ctat[3] ctl_ctat[2] ctl_ctat[1] ctl_ctat[0] start_n bandgap_core
Vdd vdd GND {vdd} 
.save v( vref )
vvref net1 vref 0
x12 vdd ptat cas net2 bandgap_cascurr_cell m=4
x13 vdd ctat cas net3 bandgap_cascurr_cell m=4
XR3 GND vref GND sky130_fd_pr__res_xhigh_po W=1 L=20 mult=1 m=1
vptat net2 net1 0
vctat net3 net1 0
Vctl_ptat4 ctl_ptat[4] GND {ctl_ptat4} 
Vctl_ptat3 ctl_ptat[3] GND {ctl_ptat3} 
Vctl_ptat2 ctl_ptat[2] GND {ctl_ptat2} 
Vctl_ptat1 ctl_ptat[1] GND {ctl_ptat1} 
Vctl_ptat0 ctl_ptat[0] GND {ctl_ptat0} 
Vctl_ctat4 ctl_ctat[4] GND {ctl_ctat4} 
Vctl_ctat3 ctl_ctat[3] GND {ctl_ctat3} 
Vctl_ctat2 ctl_ctat[2] GND {ctl_ctat2} 
Vctl_ctat1 ctl_ctat[1] GND {ctl_ctat1} 
Vctl_ctat0 ctl_ctat[0] GND {ctl_ctat0} 
Ven en GND {en} 
viout net4 net7 0
x2 vdd ptat cas net5 bandgap_cascurr_cell m=4
x3 vdd ctat cas net6 bandgap_cascurr_cell m=4
vptat2 net5 net4 0
vctat3 net6 net4 0
H1 current GND viout 1
XMmnr net7 net7 GND GND sky130_fd_pr__nfet_01v8_lvt W=1 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=3 m=3 
Vstart_n start_n GND {start_n} 
**** begin user architecture code


.temp 27
.param temp=27

*.param res_len=6.25
.param res_len=12.2

.lib sky130_fd_pr/models/sky130.lib.spice tt
.include sky130_fd_pr/models/sky130_fd_pr__model__pnp.model.spice

.param vdd=1.8

.param en=1.8
.param start_n=1.8

.param ctl_ctat4=1.8
.param ctl_ctat3=0
.param ctl_ctat2=0
.param ctl_ctat1=0
.param ctl_ctat0=0

.param ctl_ptat4=1.8
.param ctl_ptat3=0
.param ctl_ptat2=0
.param ctl_ptat1=0
.param ctl_ptat0=0

.save all
.options savecurrents

.dc temp -40 125 1


.nodeset v(xdut.q1)=1 v(xdut.q8)=1 v(xdut.ctat_r)=1

Bconverge1 xdut.q1 0 I='v(xdut.q1) < 0.0 ? 1000.0 : 0.0'
Bconverge8 xdut.q8 0 I='v(xdut.q8) < 0.0 ? 1000.0 : 0.0'
BconvergeR xdut.ctat_r 0 I='v(xdut.ctat_r) < 0.0 ? 1000.0 : 0.0'



**** end user architecture code
**.ends

* expanding   symbol:  ..//bandgap_core.sym # of pins=9

.subckt bandgap_core  vdd ptat ctat cas gnd en ctl_ptat[4] ctl_ptat[3] ctl_ptat[2] ctl_ptat[1]
+ ctl_ptat[0] ctl_ctat[4] ctl_ctat[3] ctl_ctat[2] ctl_ctat[1] ctl_ctat[0] start_n
*.iopin vdd
*.iopin gnd
*.opin ptat
*.opin ctat
*.opin cas
*.ipin en
*.ipin ctl_ptat[4],ctl_ptat[3],ctl_ptat[2],ctl_ptat[1],ctl_ptat[0]
*.ipin ctl_ctat[4],ctl_ctat[3],ctl_ctat[2],ctl_ctat[1],ctl_ctat[0]
*.ipin start_n
xop_ptat vdd ptat_int q8 q1 net15 gnd en bandgap_opamp
xop_ctat vdd ctat_int ctat_r q1 net12 gnd en bandgap_opamp
XMtri_bias_cas net1 cas vdd vdd sky130_fd_pr__pfet_01v8 W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_cas_nmirror1 net2 net2 gnd gnd sky130_fd_pr__nfet_01v8_lvt W=7 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_cas_nmirror2 cas net2 gnd gnd sky130_fd_pr__nfet_01v8_lvt W=7 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
.save v( q8 )
.save v( q8 )
.save v( ctat_r )
.save v( cas )
v2 net11 net15 0
xcurr_ptat8 vdd ptat_int cas net4 bandgap_cascurr_cell m=8
xcurr_ptat1 vdd ptat_int cas net5 bandgap_cascurr_cell m=8
xcurr_ctat vdd ctat_int cas net6 bandgap_cascurr_cell m=32
xcurr_cas_ptat vdd ptat_int cas net3 bandgap_cascurr_cell m=2
xcurr_cas_ctat vdd ctat_int cas net3 bandgap_cascurr_cell m=2
XQ1 gnd gnd q1 gnd sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ8 gnd gnd net13 gnd sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8
.save v( net11 )
xbmr net14 en bmr_biasv gnd bandgap_bmr
XMcurr_op_ptat net11 bmr_biasv vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMcurr_op_ctat net12 bmr_biasv vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMcap_ptat vdd ptat_int vdd vdd sky130_fd_pr__pfet_01v8_lvt W=7 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=32 m=32 
XMcap_ctat vdd ctat_int vdd vdd sky130_fd_pr__pfet_01v8_lvt W=7 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=64 m=64 
xtrim_ptat ctl_ptat[4] ctl_ptat[3] ctl_ptat[2] ctl_ptat[1] ctl_ptat[0] ptat net10 gnd bandgap_trim
xcurr_mirror_ptat vdd ptat_int cas net9 bandgap_cascurr_cell m=2
xtrim_ctat ctl_ctat[4] ctl_ctat[3] ctl_ctat[2] ctl_ctat[1] ctl_ctat[0] ctat net7 gnd bandgap_trim
xcurr_mirror_ctat vdd ctat_int cas net8 bandgap_cascurr_cell m=2
xcurr_ref_ptat vdd ptat cas ptat bandgap_cascurr_cell m=8
xcurr_ref_ctat vdd ctat cas ctat bandgap_cascurr_cell m=8
Vmeas1 net5 q8 0
Vmeas8 net4 q1 0
Vmeasc net6 ctat_r 0
XMsw_start q1 start_n vdd vdd sky130_fd_pr__pfet_01v8_lvt W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
Vmeas net9 net10 0
Vmeas2 net8 net7 0
.save v( bmr_biasv )
XMcas_bias cas cas net1 vdd sky130_fd_pr__pfet_01v8 W=5 L=0.5 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
Vmeas3 net3 net2 0
xres ctat_r q8 net13 gnd bandgap_resistors
XMsw_en_cas cas en vdd vdd sky130_fd_pr__pfet_01v8_hvt W=0.42 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
xen en gnd gnd vdd vdd en_n sky130_fd_sc_hd__inv_1
XMsw_en_ptatout ptat en vdd vdd sky130_fd_pr__pfet_01v8_hvt W=0.42 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en_ptatout1 ctat en vdd vdd sky130_fd_pr__pfet_01v8_hvt W=0.42 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
Vmeas4 vdd net14 0
.ends


* expanding   symbol:  bandgap_cascurr_cell/bandgap_cascurr_cell.sym # of pins=4

.subckt bandgap_cascurr_cell  vdd curr cas out
*.iopin vdd
*.ipin curr
*.ipin cas
*.opin out
XMcurr net1 curr vdd vdd sky130_fd_pr__pfet_01v8 W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMcas out cas net1 vdd sky130_fd_pr__pfet_01v8 W=5 L=0.35 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
.ends


* expanding   symbol:  bandgap_opamp/bandgap_opamp.sym # of pins=7

.subckt bandgap_opamp  vdd out inp inn bias gnd en
*.ipin inp
*.ipin inn
*.ipin bias
*.opin out
*.iopin vdd
*.iopin gnd
*.ipin en
XMcurr_diff net1 net5 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcurr_pref net5 net5 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMcurr_nref bias bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcurr_na net5 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMtriode_ncas net7 net3 gnd gnd sky130_fd_pr__nfet_01v8_lvt W=1 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_pa net3 net5 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMcas_ref net3 net3 net7 gnd sky130_fd_pr__nfet_01v8_lvt W=7 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcas_n out net3 net6 gnd sky130_fd_pr__nfet_01v8_lvt W=7 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcas_p net4 net3 net2 gnd sky130_fd_pr__nfet_01v8_lvt W=7 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcurr_loadp net4 net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_loadn out net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_foldn net6 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcurr_foldp net2 bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMdiff_n net6 inn net1 net1 sky130_fd_pr__pfet_01v8_lvt W=7 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XMdiff_p net2 inp net1 net1 sky130_fd_pr__pfet_01v8_lvt W=7 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XMsw_en_pcurr net5 en vdd vdd sky130_fd_pr__pfet_01v8_hvt W=0.42 L=8 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en_out out en_n inn gnd sky130_fd_pr__nfet_01v8 W=0.42 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en_out1 bias en_n gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
xen en gnd gnd vdd vdd en_n sky130_fd_sc_hd__inv_1
XMdumm_n gnd bias gnd gnd sky130_fd_pr__nfet_01v8_lvt W=2 L=4 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMdum_diff net1 net1 net1 net1 sky130_fd_pr__pfet_01v8_lvt W=7 L=1 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
.ends


* expanding   symbol:  bandgap_bmr/bandgap_bmr.sym # of pins=4

.subckt bandgap_bmr  vdd en biasv vss
*.iopin vdd
*.iopin vss
*.opin biasv
*.ipin en
XMdiff_n2 biasv net1 net2 vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XRbias vss net2 vss sky130_fd_pr__res_xhigh_po W=1 L=4.82 mult=1 m=1
XMdiff_n1 net1 net1 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_p2 biasv biasv vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMcurr_p1 net1 biasv vdd vdd sky130_fd_pr__pfet_01v8_lvt W=5 L=8 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_start net5 net3 net1 vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMdiff_n3 net3 net1 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_bias net3 net3 vdd vdd sky130_fd_pr__pfet_01v8_lvt W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)'
+ as='W * 0.29' ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en_p biasv en vdd vdd sky130_fd_pr__pfet_01v8 W=0.42 L=4.00 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XCcomp biasv net1 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
XMdum2 vss net1 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XCfilt biasv vdd sky130_fd_pr__cap_mim_m3_1 W=7.2 L=7.7 MF=1 m=1
XMdum1 vss net3 vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_en_n net1 net4 vss vss sky130_fd_pr__nfet_01v8 W=0.42 L=1.00 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
xen en vss vss vdd vdd net4 sky130_fd_sc_hd__inv_1
XMsw_en_n1 biasv en net5 vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMdum3 vss en vss vss sky130_fd_pr__nfet_01v8 W=5 L=1 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
.ends


* expanding   symbol:  bandgap_trim/bandgap_trim.sym # of pins=4

.subckt bandgap_trim  ctl[4] ctl[3] ctl[2] ctl[1] ctl[0] out in gnd
*.ipin ctl[4],ctl[3],ctl[2],ctl[1],ctl[0]
*.ipin gnd
*.ipin in
*.opin out
XMcurr_3 net2 in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMcurr_2 net3 in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMcurr_1 net4 in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMcurr_0 net5 in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMsw_3 out ctl[3] net2 gnd sky130_fd_pr__nfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=8 m=8 
XMsw_2 out ctl[2] net3 gnd sky130_fd_pr__nfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=4 m=4 
XMsw_1 out ctl[1] net4 gnd sky130_fd_pr__nfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=2 m=2 
XMsw_0 out ctl[0] net5 gnd sky130_fd_pr__nfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=1 m=1 
XMcurr_4 net1 in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XMsw_4 out ctl[4] net1 gnd sky130_fd_pr__nfet_01v8 W=0.42 L=0.15 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XMcurr_ref in in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=16 m=16 
XMcurr_base out in gnd gnd sky130_fd_pr__nfet_01v8 W=0.42 L=20 ad='W * 0.29' pd='2 * (W + 0.29)' as='W * 0.29'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 nf=1 mult=48 m=48 
.ends


* expanding   symbol:  bandgap_resistors/bandgap_resistors.sym # of pins=4

.subckt bandgap_resistors  ctat ptat1 ptat2 gnd
*.iopin ptat1
*.iopin ptat2
*.iopin gnd
*.iopin ctat
XRptat3 ptat2 net1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat5 ptat2 net1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat2 net1 ptat1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat1 net1 ptat1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat8 ptat2 net1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat7 ptat2 net1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat4 net1 ptat1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRptat6 net1 ptat1 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat2 net2 ctat gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat1 net2 ctat gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat6 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat5 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat8 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat7 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat9 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat11 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat10 gnd net3 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat3 net3 net2 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRctat4 net3 net2 gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRdumm2 gnd gnd gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
XRdumm1 gnd gnd gnd sky130_fd_pr__res_xhigh_po W=1 L=12.4 mult=1 m=1
.ends

.GLOBAL GND
**** begin user architecture code
.include /home/tom/repositories/amsat_txrx_ic/../skywater/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_1.spice

**** end user architecture code
.end
